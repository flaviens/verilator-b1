// Copyright 2023 Flavien Solt, ETH Zurich.
// Licensed under the General Public License, Version 3.0, see LICENSE for details.
// SPDX-License-Identifier: GPL-3.0-only

module top(in_data, out_data);
  input [262143:0] in_data;
  wire [262143:0] in_data;
  output [131071:0] out_data;
  wire [131071:0] out_data;
  assign out_data[799:768] = in_data[1567:1536] - in_data[1599:1568];
  assign out_data[7999:7968] = in_data[15967:15936] - in_data[15999:15968];
  assign out_data[79999:79968] = in_data[159967:159936] - in_data[159999:159968];
  assign out_data[80031:80000] = in_data[160031:160000] - in_data[160063:160032];
  assign out_data[80063:80032] = in_data[160095:160064] - in_data[160127:160096];
  assign out_data[80095:80064] = in_data[160159:160128] - in_data[160191:160160];
  assign out_data[80127:80096] = in_data[160223:160192] - in_data[160255:160224];
  assign out_data[80159:80128] = in_data[160287:160256] - in_data[160319:160288];
  assign out_data[80191:80160] = in_data[160351:160320] - in_data[160383:160352];
  assign out_data[80223:80192] = in_data[160415:160384] - in_data[160447:160416];
  assign out_data[80255:80224] = in_data[160479:160448] - in_data[160511:160480];
  assign out_data[80287:80256] = in_data[160543:160512] - in_data[160575:160544];
  assign out_data[8031:8000] = in_data[16031:16000] - in_data[16063:16032];
  assign out_data[80351:80320] = in_data[160671:160640] - in_data[160703:160672];
  assign out_data[80383:80352] = in_data[160735:160704] - in_data[160767:160736];
  assign out_data[80415:80384] = in_data[160799:160768] - in_data[160831:160800];
  assign out_data[80447:80416] = in_data[160863:160832] - in_data[160895:160864];
  assign out_data[80479:80448] = in_data[160927:160896] - in_data[160959:160928];
  assign out_data[80511:80480] = in_data[160991:160960] - in_data[161023:160992];
  assign out_data[80543:80512] = in_data[161055:161024] - in_data[161087:161056];
  assign out_data[80575:80544] = in_data[161119:161088] - in_data[161151:161120];
  assign out_data[80607:80576] = in_data[161183:161152] - in_data[161215:161184];
  assign out_data[8063:8032] = in_data[16095:16064] - in_data[16127:16096];
  assign out_data[80639:80608] = in_data[161247:161216] - in_data[161279:161248];
  assign out_data[80671:80640] = in_data[161311:161280] - in_data[161343:161312];
  assign out_data[80799:80768] = in_data[161567:161536] - in_data[161599:161568];
  assign out_data[80831:80800] = in_data[161631:161600] - in_data[161663:161632];
  assign out_data[80863:80832] = in_data[161695:161664] - in_data[161727:161696];
  assign out_data[80895:80864] = in_data[161759:161728] - in_data[161791:161760];
  assign out_data[80927:80896] = in_data[161823:161792] - in_data[161855:161824];
  assign out_data[8095:8064] = in_data[16159:16128] - in_data[16191:16160];
  assign out_data[80959:80928] = in_data[161887:161856] - in_data[161919:161888];
  assign out_data[80991:80960] = in_data[161951:161920] - in_data[161983:161952];
  assign out_data[81023:80992] = in_data[162015:161984] - in_data[162047:162016];
  assign out_data[81055:81024] = in_data[162079:162048] - in_data[162111:162080];
  assign out_data[81087:81056] = in_data[162143:162112] - in_data[162175:162144];
  assign out_data[81119:81088] = in_data[162207:162176] - in_data[162239:162208];
  assign out_data[81151:81120] = in_data[162271:162240] - in_data[162303:162272];
  assign out_data[81183:81152] = in_data[162335:162304] - in_data[162367:162336];
  assign out_data[81215:81184] = in_data[162399:162368] - in_data[162431:162400];
  assign out_data[81247:81216] = in_data[162463:162432] - in_data[162495:162464];
  assign out_data[8127:8096] = in_data[16223:16192] - in_data[16255:16224];
  assign out_data[81279:81248] = in_data[162527:162496] - in_data[162559:162528];
  assign out_data[81311:81280] = in_data[162591:162560] - in_data[162623:162592];
  assign out_data[81343:81312] = in_data[162655:162624] - in_data[162687:162656];
  assign out_data[81375:81344] = in_data[162719:162688] - in_data[162751:162720];
  assign out_data[81407:81376] = in_data[162783:162752] - in_data[162815:162784];
  assign out_data[81439:81408] = in_data[162847:162816] - in_data[162879:162848];
  assign out_data[81471:81440] = in_data[162911:162880] - in_data[162943:162912];
  assign out_data[81503:81472] = in_data[162975:162944] - in_data[163007:162976];
  assign out_data[81535:81504] = in_data[163039:163008] - in_data[163071:163040];
  assign out_data[81567:81536] = in_data[163103:163072] - in_data[163135:163104];
  assign out_data[8159:8128] = in_data[16287:16256] - in_data[16319:16288];
  assign out_data[81599:81568] = in_data[163167:163136] - in_data[163199:163168];
  assign out_data[81631:81600] = in_data[163231:163200] - in_data[163263:163232];
  assign out_data[81663:81632] = in_data[163295:163264] - in_data[163327:163296];
  assign out_data[81695:81664] = in_data[163359:163328] - in_data[163391:163360];
  assign out_data[81727:81696] = in_data[163423:163392] - in_data[163455:163424];
  assign out_data[81759:81728] = in_data[163487:163456] - in_data[163519:163488];
  assign out_data[81791:81760] = in_data[163551:163520] - in_data[163583:163552];
  assign out_data[81823:81792] = in_data[163615:163584] - in_data[163647:163616];
  assign out_data[81855:81824] = in_data[163679:163648] - in_data[163711:163680];
  assign out_data[81887:81856] = in_data[163743:163712] - in_data[163775:163744];
  assign out_data[8191:8160] = in_data[16351:16320] - in_data[16383:16352];
  assign out_data[81919:81888] = in_data[163807:163776] - in_data[163839:163808];
  assign out_data[81951:81920] = in_data[163871:163840] - in_data[163903:163872];
  assign out_data[81983:81952] = in_data[163935:163904] - in_data[163967:163936];
  assign out_data[82015:81984] = in_data[163999:163968] - in_data[164031:164000];
  assign out_data[82047:82016] = in_data[164063:164032] - in_data[164095:164064];
  assign out_data[82079:82048] = in_data[164127:164096] - in_data[164159:164128];
  assign out_data[82111:82080] = in_data[164191:164160] - in_data[164223:164192];
  assign out_data[82143:82112] = in_data[164255:164224] - in_data[164287:164256];
  assign out_data[82175:82144] = in_data[164319:164288] - in_data[164351:164320];
  assign out_data[82207:82176] = in_data[164383:164352] - in_data[164415:164384];
  assign out_data[8223:8192] = in_data[16415:16384] - in_data[16447:16416];
  assign out_data[82239:82208] = in_data[164447:164416] - in_data[164479:164448];
  assign out_data[82271:82240] = in_data[164511:164480] - in_data[164543:164512];
  assign out_data[82303:82272] = in_data[164575:164544] - in_data[164607:164576];
  assign out_data[82335:82304] = in_data[164639:164608] - in_data[164671:164640];
  assign out_data[82367:82336] = in_data[164703:164672] - in_data[164735:164704];
  assign out_data[82399:82368] = in_data[164767:164736] - in_data[164799:164768];
  assign out_data[82431:82400] = in_data[164831:164800] - in_data[164863:164832];
  assign out_data[82463:82432] = in_data[164895:164864] - in_data[164927:164896];
  assign out_data[82495:82464] = in_data[164959:164928] - in_data[164991:164960];
  assign out_data[82527:82496] = in_data[165023:164992] - in_data[165055:165024];
  assign out_data[8255:8224] = in_data[16479:16448] - in_data[16511:16480];
  assign out_data[82559:82528] = in_data[165087:165056] - in_data[165119:165088];
  assign out_data[82591:82560] = in_data[165151:165120] - in_data[165183:165152];
  assign out_data[82623:82592] = in_data[165215:165184] - in_data[165247:165216];
  assign out_data[82655:82624] = in_data[165279:165248] - in_data[165311:165280];
  assign out_data[82687:82656] = in_data[165343:165312] - in_data[165375:165344];
  assign out_data[82719:82688] = in_data[165407:165376] - in_data[165439:165408];
  assign out_data[82751:82720] = in_data[165471:165440] - in_data[165503:165472];
  assign out_data[82783:82752] = in_data[165535:165504] - in_data[165567:165536];
  assign out_data[82815:82784] = in_data[165599:165568] - in_data[165631:165600];
  assign out_data[82847:82816] = in_data[165663:165632] - in_data[165695:165664];
  assign out_data[8287:8256] = in_data[16543:16512] - in_data[16575:16544];
  assign out_data[82879:82848] = in_data[165727:165696] - in_data[165759:165728];
  assign out_data[82911:82880] = in_data[165791:165760] - in_data[165823:165792];
  assign out_data[82943:82912] = in_data[165855:165824] - in_data[165887:165856];
  assign out_data[82975:82944] = in_data[165919:165888] - in_data[165951:165920];
  assign out_data[83007:82976] = in_data[165983:165952] - in_data[166015:165984];
  assign out_data[83039:83008] = in_data[166047:166016] - in_data[166079:166048];
  assign out_data[83071:83040] = in_data[166111:166080] - in_data[166143:166112];
  assign out_data[83103:83072] = in_data[166175:166144] - in_data[166207:166176];
  assign out_data[83135:83104] = in_data[166239:166208] - in_data[166271:166240];
  assign out_data[83167:83136] = in_data[166303:166272] - in_data[166335:166304];
  assign out_data[831:800] = in_data[1631:1600] - in_data[1663:1632];
  assign out_data[8319:8288] = in_data[16607:16576] - in_data[16639:16608];
  assign out_data[83199:83168] = in_data[166367:166336] - in_data[166399:166368];
  assign out_data[83231:83200] = in_data[166431:166400] - in_data[166463:166432];
  assign out_data[83263:83232] = in_data[166495:166464] - in_data[166527:166496];
  assign out_data[83295:83264] = in_data[166559:166528] - in_data[166591:166560];
  assign out_data[83327:83296] = in_data[166623:166592] - in_data[166655:166624];
  assign out_data[83359:83328] = in_data[166687:166656] - in_data[166719:166688];
  assign out_data[83391:83360] = in_data[166751:166720] - in_data[166783:166752];
  assign out_data[83423:83392] = in_data[166815:166784] - in_data[166847:166816];
  assign out_data[83455:83424] = in_data[166879:166848] - in_data[166911:166880];
  assign out_data[83487:83456] = in_data[166943:166912] - in_data[166975:166944];
  assign out_data[8351:8320] = in_data[16671:16640] - in_data[16703:16672];
  assign out_data[83519:83488] = in_data[167007:166976] - in_data[167039:167008];
  assign out_data[83551:83520] = in_data[167071:167040] - in_data[167103:167072];
  assign out_data[83583:83552] = in_data[167135:167104] - in_data[167167:167136];
  assign out_data[83615:83584] = in_data[167199:167168] - in_data[167231:167200];
  assign out_data[83647:83616] = in_data[167263:167232] - in_data[167295:167264];
  assign out_data[83679:83648] = in_data[167327:167296] - in_data[167359:167328];
  assign out_data[83711:83680] = in_data[167391:167360] - in_data[167423:167392];
  assign out_data[83743:83712] = in_data[167455:167424] - in_data[167487:167456];
  assign out_data[83775:83744] = in_data[167519:167488] - in_data[167551:167520];
  assign out_data[83807:83776] = in_data[167583:167552] - in_data[167615:167584];
  assign out_data[8383:8352] = in_data[16735:16704] - in_data[16767:16736];
  assign out_data[83839:83808] = in_data[167647:167616] - in_data[167679:167648];
  assign out_data[83871:83840] = in_data[167711:167680] - in_data[167743:167712];
  assign out_data[83903:83872] = in_data[167775:167744] - in_data[167807:167776];
  assign out_data[83935:83904] = in_data[167839:167808] - in_data[167871:167840];
  assign out_data[83967:83936] = in_data[167903:167872] - in_data[167935:167904];
  assign out_data[83999:83968] = in_data[167967:167936] - in_data[167999:167968];
  assign out_data[84031:84000] = in_data[168031:168000] - in_data[168063:168032];
  assign out_data[84063:84032] = in_data[168095:168064] - in_data[168127:168096];
  assign out_data[84095:84064] = in_data[168159:168128] - in_data[168191:168160];
  assign out_data[84127:84096] = in_data[168223:168192] - in_data[168255:168224];
  assign out_data[8415:8384] = in_data[16799:16768] - in_data[16831:16800];
  assign out_data[84159:84128] = in_data[168287:168256] - in_data[168319:168288];
  assign out_data[84191:84160] = in_data[168351:168320] - in_data[168383:168352];
  assign out_data[84223:84192] = in_data[168415:168384] - in_data[168447:168416];
  assign out_data[84255:84224] = in_data[168479:168448] - in_data[168511:168480];
  assign out_data[84287:84256] = in_data[168543:168512] - in_data[168575:168544];
  assign out_data[84319:84288] = in_data[168607:168576] - in_data[168639:168608];
  assign out_data[84351:84320] = in_data[168671:168640] - in_data[168703:168672];
  assign out_data[84383:84352] = in_data[168735:168704] - in_data[168767:168736];
  assign out_data[84415:84384] = in_data[168799:168768] - in_data[168831:168800];
  assign out_data[84447:84416] = in_data[168863:168832] - in_data[168895:168864];
  assign out_data[8447:8416] = in_data[16863:16832] - in_data[16895:16864];
  assign out_data[84479:84448] = in_data[168927:168896] - in_data[168959:168928];
  assign out_data[84511:84480] = in_data[168991:168960] - in_data[169023:168992];
  assign out_data[84543:84512] = in_data[169055:169024] - in_data[169087:169056];
  assign out_data[84575:84544] = in_data[169119:169088] - in_data[169151:169120];
  assign out_data[84607:84576] = in_data[169183:169152] - in_data[169215:169184];
  assign out_data[84639:84608] = in_data[169247:169216] - in_data[169279:169248];
  assign out_data[84671:84640] = in_data[169311:169280] - in_data[169343:169312];
  assign out_data[84703:84672] = in_data[169375:169344] - in_data[169407:169376];
  assign out_data[84735:84704] = in_data[169439:169408] - in_data[169471:169440];
  assign out_data[84767:84736] = in_data[169503:169472] - in_data[169535:169504];
  assign out_data[8479:8448] = in_data[16927:16896] - in_data[16959:16928];
  assign out_data[84799:84768] = in_data[169567:169536] - in_data[169599:169568];
  assign out_data[84831:84800] = in_data[169631:169600] - in_data[169663:169632];
  assign out_data[84863:84832] = in_data[169695:169664] - in_data[169727:169696];
  assign out_data[84895:84864] = in_data[169759:169728] - in_data[169791:169760];
  assign out_data[84927:84896] = in_data[169823:169792] - in_data[169855:169824];
  assign out_data[84959:84928] = in_data[169887:169856] - in_data[169919:169888];
  assign out_data[84991:84960] = in_data[169951:169920] - in_data[169983:169952];
  assign out_data[85023:84992] = in_data[170015:169984] - in_data[170047:170016];
  assign out_data[85055:85024] = in_data[170079:170048] - in_data[170111:170080];
  assign out_data[85087:85056] = in_data[170143:170112] - in_data[170175:170144];
  assign out_data[8511:8480] = in_data[16991:16960] - in_data[17023:16992];
  assign out_data[85119:85088] = in_data[170207:170176] - in_data[170239:170208];
  assign out_data[85151:85120] = in_data[170271:170240] - in_data[170303:170272];
  assign out_data[85183:85152] = in_data[170335:170304] - in_data[170367:170336];
  assign out_data[85215:85184] = in_data[170399:170368] - in_data[170431:170400];
  assign out_data[85247:85216] = in_data[170463:170432] - in_data[170495:170464];
  assign out_data[85279:85248] = in_data[170527:170496] - in_data[170559:170528];
  assign out_data[85311:85280] = in_data[170591:170560] - in_data[170623:170592];
  assign out_data[85343:85312] = in_data[170655:170624] - in_data[170687:170656];
  assign out_data[85375:85344] = in_data[170719:170688] - in_data[170751:170720];
  assign out_data[85407:85376] = in_data[170783:170752] - in_data[170815:170784];
  assign out_data[8543:8512] = in_data[17055:17024] - in_data[17087:17056];
  assign out_data[85439:85408] = in_data[170847:170816] - in_data[170879:170848];
  assign out_data[85471:85440] = in_data[170911:170880] - in_data[170943:170912];
  assign out_data[85503:85472] = in_data[170975:170944] - in_data[171007:170976];
  assign out_data[85535:85504] = in_data[171039:171008] - in_data[171071:171040];
  assign out_data[85567:85536] = in_data[171103:171072] - in_data[171135:171104];
  assign out_data[85599:85568] = in_data[171167:171136] - in_data[171199:171168];
  assign out_data[85631:85600] = in_data[171231:171200] - in_data[171263:171232];
  assign out_data[85663:85632] = in_data[171295:171264] - in_data[171327:171296];
  assign out_data[85695:85664] = in_data[171359:171328] - in_data[171391:171360];
  assign out_data[85727:85696] = in_data[171423:171392] - in_data[171455:171424];
  assign out_data[8575:8544] = in_data[17119:17088] - in_data[17151:17120];
  assign out_data[85759:85728] = in_data[171487:171456] - in_data[171519:171488];
  assign out_data[85791:85760] = in_data[171551:171520] - in_data[171583:171552];
  assign out_data[85823:85792] = in_data[171615:171584] - in_data[171647:171616];
  assign out_data[85855:85824] = in_data[171679:171648] - in_data[171711:171680];
  assign out_data[85887:85856] = in_data[171743:171712] - in_data[171775:171744];
  assign out_data[85919:85888] = in_data[171807:171776] - in_data[171839:171808];
  assign out_data[85951:85920] = in_data[171871:171840] - in_data[171903:171872];
  assign out_data[85983:85952] = in_data[171935:171904] - in_data[171967:171936];
  assign out_data[86015:85984] = in_data[171999:171968] - in_data[172031:172000];
  assign out_data[86047:86016] = in_data[172063:172032] - in_data[172095:172064];
  assign out_data[8607:8576] = in_data[17183:17152] - in_data[17215:17184];
  assign out_data[86079:86048] = in_data[172127:172096] - in_data[172159:172128];
  assign out_data[86111:86080] = in_data[172191:172160] - in_data[172223:172192];
  assign out_data[86143:86112] = in_data[172255:172224] - in_data[172287:172256];
  assign out_data[86175:86144] = in_data[172319:172288] - in_data[172351:172320];
  assign out_data[86207:86176] = in_data[172383:172352] - in_data[172415:172384];
  assign out_data[86239:86208] = in_data[172447:172416] - in_data[172479:172448];
  assign out_data[86271:86240] = in_data[172511:172480] - in_data[172543:172512];
  assign out_data[86303:86272] = in_data[172575:172544] - in_data[172607:172576];
  assign out_data[86335:86304] = in_data[172639:172608] - in_data[172671:172640];
  assign out_data[86367:86336] = in_data[172703:172672] - in_data[172735:172704];
  assign out_data[863:832] = in_data[1695:1664] - in_data[1727:1696];
  assign out_data[8639:8608] = in_data[17247:17216] - in_data[17279:17248];
  assign out_data[86399:86368] = in_data[172767:172736] - in_data[172799:172768];
  assign out_data[86431:86400] = in_data[172831:172800] - in_data[172863:172832];
  assign out_data[86463:86432] = in_data[172895:172864] - in_data[172927:172896];
  assign out_data[86495:86464] = in_data[172959:172928] - in_data[172991:172960];
  assign out_data[86527:86496] = in_data[173023:172992] - in_data[173055:173024];
  assign out_data[86559:86528] = in_data[173087:173056] - in_data[173119:173088];
  assign out_data[86591:86560] = in_data[173151:173120] - in_data[173183:173152];
  assign out_data[86623:86592] = in_data[173215:173184] - in_data[173247:173216];
  assign out_data[86655:86624] = in_data[173279:173248] - in_data[173311:173280];
  assign out_data[86687:86656] = in_data[173343:173312] - in_data[173375:173344];
  assign out_data[8671:8640] = in_data[17311:17280] - in_data[17343:17312];
  assign out_data[86719:86688] = in_data[173407:173376] - in_data[173439:173408];
  assign out_data[86751:86720] = in_data[173471:173440] - in_data[173503:173472];
  assign out_data[86783:86752] = in_data[173535:173504] - in_data[173567:173536];
  assign out_data[86815:86784] = in_data[173599:173568] - in_data[173631:173600];
  assign out_data[86847:86816] = in_data[173663:173632] - in_data[173695:173664];
  assign out_data[86879:86848] = in_data[173727:173696] - in_data[173759:173728];
  assign out_data[86911:86880] = in_data[173791:173760] - in_data[173823:173792];
  assign out_data[86943:86912] = in_data[173855:173824] - in_data[173887:173856];
  assign out_data[86975:86944] = in_data[173919:173888] - in_data[173951:173920];
  assign out_data[87007:86976] = in_data[173983:173952] - in_data[174015:173984];
  assign out_data[8703:8672] = in_data[17375:17344] - in_data[17407:17376];
  assign out_data[87039:87008] = in_data[174047:174016] - in_data[174079:174048];
  assign out_data[87071:87040] = in_data[174111:174080] - in_data[174143:174112];
  assign out_data[87103:87072] = in_data[174175:174144] - in_data[174207:174176];
  assign out_data[87135:87104] = in_data[174239:174208] - in_data[174271:174240];
  assign out_data[87167:87136] = in_data[174303:174272] - in_data[174335:174304];
  assign out_data[87199:87168] = in_data[174367:174336] - in_data[174399:174368];
  assign out_data[87231:87200] = in_data[174431:174400] - in_data[174463:174432];
  assign out_data[87263:87232] = in_data[174495:174464] - in_data[174527:174496];
  assign out_data[87295:87264] = in_data[174559:174528] - in_data[174591:174560];
  assign out_data[87327:87296] = in_data[174623:174592] - in_data[174655:174624];
  assign out_data[8735:8704] = in_data[17439:17408] - in_data[17471:17440];
  assign out_data[87359:87328] = in_data[174687:174656] - in_data[174719:174688];
  assign out_data[87391:87360] = in_data[174751:174720] - in_data[174783:174752];
  assign out_data[87423:87392] = in_data[174815:174784] - in_data[174847:174816];
  assign out_data[87455:87424] = in_data[174879:174848] - in_data[174911:174880];
  assign out_data[87487:87456] = in_data[174943:174912] - in_data[174975:174944];
  assign out_data[87519:87488] = in_data[175007:174976] - in_data[175039:175008];
  assign out_data[87551:87520] = in_data[175071:175040] - in_data[175103:175072];
  assign out_data[87583:87552] = in_data[175135:175104] - in_data[175167:175136];
  assign out_data[87615:87584] = in_data[175199:175168] - in_data[175231:175200];
  assign out_data[87647:87616] = in_data[175263:175232] - in_data[175295:175264];
  assign out_data[8767:8736] = in_data[17503:17472] - in_data[17535:17504];
  assign out_data[87679:87648] = in_data[175327:175296] - in_data[175359:175328];
  assign out_data[87711:87680] = in_data[175391:175360] - in_data[175423:175392];
  assign out_data[87743:87712] = in_data[175455:175424] - in_data[175487:175456];
  assign out_data[87775:87744] = in_data[175519:175488] - in_data[175551:175520];
  assign out_data[87807:87776] = in_data[175583:175552] - in_data[175615:175584];
  assign out_data[87839:87808] = in_data[175647:175616] - in_data[175679:175648];
  assign out_data[87871:87840] = in_data[175711:175680] - in_data[175743:175712];
  assign out_data[87903:87872] = in_data[175775:175744] - in_data[175807:175776];
  assign out_data[87935:87904] = in_data[175839:175808] - in_data[175871:175840];
  assign out_data[87967:87936] = in_data[175903:175872] - in_data[175935:175904];
  assign out_data[8799:8768] = in_data[17567:17536] - in_data[17599:17568];
  assign out_data[87999:87968] = in_data[175967:175936] - in_data[175999:175968];
  assign out_data[88031:88000] = in_data[176031:176000] - in_data[176063:176032];
  assign out_data[88063:88032] = in_data[176095:176064] - in_data[176127:176096];
  assign out_data[88095:88064] = in_data[176159:176128] - in_data[176191:176160];
  assign out_data[88127:88096] = in_data[176223:176192] - in_data[176255:176224];
  assign out_data[88159:88128] = in_data[176287:176256] - in_data[176319:176288];
  assign out_data[88191:88160] = in_data[176351:176320] - in_data[176383:176352];
  assign out_data[88223:88192] = in_data[176415:176384] - in_data[176447:176416];
  assign out_data[88255:88224] = in_data[176479:176448] - in_data[176511:176480];
  assign out_data[88287:88256] = in_data[176543:176512] - in_data[176575:176544];
  assign out_data[8831:8800] = in_data[17631:17600] - in_data[17663:17632];
  assign out_data[88319:88288] = in_data[176607:176576] - in_data[176639:176608];
  assign out_data[88351:88320] = in_data[176671:176640] - in_data[176703:176672];
  assign out_data[88383:88352] = in_data[176735:176704] - in_data[176767:176736];
  assign out_data[88415:88384] = in_data[176799:176768] - in_data[176831:176800];
  assign out_data[88447:88416] = in_data[176863:176832] - in_data[176895:176864];
  assign out_data[88479:88448] = in_data[176927:176896] - in_data[176959:176928];
  assign out_data[88511:88480] = in_data[176991:176960] - in_data[177023:176992];
  assign out_data[88543:88512] = in_data[177055:177024] - in_data[177087:177056];
  assign out_data[88575:88544] = in_data[177119:177088] - in_data[177151:177120];
  assign out_data[88607:88576] = in_data[177183:177152] - in_data[177215:177184];
  assign out_data[8863:8832] = in_data[17695:17664] - in_data[17727:17696];
  assign out_data[88639:88608] = in_data[177247:177216] - in_data[177279:177248];
  assign out_data[88671:88640] = in_data[177311:177280] - in_data[177343:177312];
  assign out_data[88703:88672] = in_data[177375:177344] - in_data[177407:177376];
  assign out_data[88735:88704] = in_data[177439:177408] - in_data[177471:177440];
  assign out_data[88767:88736] = in_data[177503:177472] - in_data[177535:177504];
  assign out_data[88799:88768] = in_data[177567:177536] - in_data[177599:177568];
  assign out_data[88831:88800] = in_data[177631:177600] - in_data[177663:177632];
  assign out_data[88863:88832] = in_data[177695:177664] - in_data[177727:177696];
  assign out_data[88895:88864] = in_data[177759:177728] - in_data[177791:177760];
  assign out_data[88927:88896] = in_data[177823:177792] - in_data[177855:177824];
  assign out_data[8895:8864] = in_data[17759:17728] - in_data[17791:17760];
  assign out_data[88959:88928] = in_data[177887:177856] - in_data[177919:177888];
  assign out_data[88991:88960] = in_data[177951:177920] - in_data[177983:177952];
  assign out_data[89023:88992] = in_data[178015:177984] - in_data[178047:178016];
  assign out_data[89055:89024] = in_data[178079:178048] - in_data[178111:178080];
  assign out_data[89087:89056] = in_data[178143:178112] - in_data[178175:178144];
  assign out_data[89119:89088] = in_data[178207:178176] - in_data[178239:178208];
  assign out_data[89151:89120] = in_data[178271:178240] - in_data[178303:178272];
  assign out_data[89183:89152] = in_data[178335:178304] - in_data[178367:178336];
  assign out_data[89215:89184] = in_data[178399:178368] - in_data[178431:178400];
  assign out_data[89247:89216] = in_data[178463:178432] - in_data[178495:178464];
  assign out_data[8927:8896] = in_data[17823:17792] - in_data[17855:17824];
  assign out_data[89279:89248] = in_data[178527:178496] - in_data[178559:178528];
  assign out_data[89311:89280] = in_data[178591:178560] - in_data[178623:178592];
  assign out_data[89343:89312] = in_data[178655:178624] - in_data[178687:178656];
  assign out_data[89375:89344] = in_data[178719:178688] - in_data[178751:178720];
  assign out_data[89407:89376] = in_data[178783:178752] - in_data[178815:178784];
  assign out_data[89439:89408] = in_data[178847:178816] - in_data[178879:178848];
  assign out_data[89471:89440] = in_data[178911:178880] - in_data[178943:178912];
  assign out_data[89503:89472] = in_data[178975:178944] - in_data[179007:178976];
  assign out_data[89535:89504] = in_data[179039:179008] - in_data[179071:179040];
  assign out_data[89567:89536] = in_data[179103:179072] - in_data[179135:179104];
  assign out_data[895:864] = in_data[1759:1728] - in_data[1791:1760];
  assign out_data[8959:8928] = in_data[17887:17856] - in_data[17919:17888];
  assign out_data[89599:89568] = in_data[179167:179136] - in_data[179199:179168];
  assign out_data[89631:89600] = in_data[179231:179200] - in_data[179263:179232];
  assign out_data[89663:89632] = in_data[179295:179264] - in_data[179327:179296];
  assign out_data[89695:89664] = in_data[179359:179328] - in_data[179391:179360];
  assign out_data[89727:89696] = in_data[179423:179392] - in_data[179455:179424];
  assign out_data[89759:89728] = in_data[179487:179456] - in_data[179519:179488];
  assign out_data[89791:89760] = in_data[179551:179520] - in_data[179583:179552];
  assign out_data[89823:89792] = in_data[179615:179584] - in_data[179647:179616];
  assign out_data[89855:89824] = in_data[179679:179648] - in_data[179711:179680];
  assign out_data[89887:89856] = in_data[179743:179712] - in_data[179775:179744];
  assign out_data[8991:8960] = in_data[17951:17920] - in_data[17983:17952];
  assign out_data[89919:89888] = in_data[179807:179776] - in_data[179839:179808];
  assign out_data[89951:89920] = in_data[179871:179840] - in_data[179903:179872];
  assign out_data[89983:89952] = in_data[179935:179904] - in_data[179967:179936];
  assign out_data[90015:89984] = in_data[179999:179968] - in_data[180031:180000];
  assign out_data[90047:90016] = in_data[180063:180032] - in_data[180095:180064];
  assign out_data[90079:90048] = in_data[180127:180096] - in_data[180159:180128];
  assign out_data[90111:90080] = in_data[180191:180160] - in_data[180223:180192];
  assign out_data[90143:90112] = in_data[180255:180224] - in_data[180287:180256];
  assign out_data[90175:90144] = in_data[180319:180288] - in_data[180351:180320];
  assign out_data[90207:90176] = in_data[180383:180352] - in_data[180415:180384];
  assign out_data[9023:8992] = in_data[18015:17984] - in_data[18047:18016];
  assign out_data[90239:90208] = in_data[180447:180416] - in_data[180479:180448];
  assign out_data[90271:90240] = in_data[180511:180480] - in_data[180543:180512];
  assign out_data[90303:90272] = in_data[180575:180544] - in_data[180607:180576];
  assign out_data[90335:90304] = in_data[180639:180608] - in_data[180671:180640];
  assign out_data[90367:90336] = in_data[180703:180672] - in_data[180735:180704];
  assign out_data[90399:90368] = in_data[180767:180736] - in_data[180799:180768];
  assign out_data[90431:90400] = in_data[180831:180800] - in_data[180863:180832];
  assign out_data[90463:90432] = in_data[180895:180864] - in_data[180927:180896];
  assign out_data[90495:90464] = in_data[180959:180928] - in_data[180991:180960];
  assign out_data[90527:90496] = in_data[181023:180992] - in_data[181055:181024];
  assign out_data[9055:9024] = in_data[18079:18048] - in_data[18111:18080];
  assign out_data[90559:90528] = in_data[181087:181056] - in_data[181119:181088];
  assign out_data[90591:90560] = in_data[181151:181120] - in_data[181183:181152];
  assign out_data[90623:90592] = in_data[181215:181184] - in_data[181247:181216];
  assign out_data[90655:90624] = in_data[181279:181248] - in_data[181311:181280];
  assign out_data[90687:90656] = in_data[181343:181312] - in_data[181375:181344];
  assign out_data[90719:90688] = in_data[181407:181376] - in_data[181439:181408];
  assign out_data[90751:90720] = in_data[181471:181440] - in_data[181503:181472];
  assign out_data[90783:90752] = in_data[181535:181504] - in_data[181567:181536];
  assign out_data[90815:90784] = in_data[181599:181568] - in_data[181631:181600];
  assign out_data[90847:90816] = in_data[181663:181632] - in_data[181695:181664];
  assign out_data[9087:9056] = in_data[18143:18112] - in_data[18175:18144];
  assign out_data[90879:90848] = in_data[181727:181696] - in_data[181759:181728];
  assign out_data[90911:90880] = in_data[181791:181760] - in_data[181823:181792];
  assign out_data[90943:90912] = in_data[181855:181824] - in_data[181887:181856];
  assign out_data[90975:90944] = in_data[181919:181888] - in_data[181951:181920];
  assign out_data[91007:90976] = in_data[181983:181952] - in_data[182015:181984];
  assign out_data[91039:91008] = in_data[182047:182016] - in_data[182079:182048];
  assign out_data[91071:91040] = in_data[182111:182080] - in_data[182143:182112];
  assign out_data[91103:91072] = in_data[182175:182144] - in_data[182207:182176];
  assign out_data[91135:91104] = in_data[182239:182208] - in_data[182271:182240];
  assign out_data[91167:91136] = in_data[182303:182272] - in_data[182335:182304];
  assign out_data[9119:9088] = in_data[18207:18176] - in_data[18239:18208];
  assign out_data[91199:91168] = in_data[182367:182336] - in_data[182399:182368];
  assign out_data[91231:91200] = in_data[182431:182400] - in_data[182463:182432];
  assign out_data[91263:91232] = in_data[182495:182464] - in_data[182527:182496];
  assign out_data[91295:91264] = in_data[182559:182528] - in_data[182591:182560];
  assign out_data[91327:91296] = in_data[182623:182592] - in_data[182655:182624];
  assign out_data[91359:91328] = in_data[182687:182656] - in_data[182719:182688];
  assign out_data[91391:91360] = in_data[182751:182720] - in_data[182783:182752];
  assign out_data[91423:91392] = in_data[182815:182784] - in_data[182847:182816];
  assign out_data[91455:91424] = in_data[182879:182848] - in_data[182911:182880];
  assign out_data[91487:91456] = in_data[182943:182912] - in_data[182975:182944];
  assign out_data[9151:9120] = in_data[18271:18240] - in_data[18303:18272];
  assign out_data[91519:91488] = in_data[183007:182976] - in_data[183039:183008];
  assign out_data[91551:91520] = in_data[183071:183040] - in_data[183103:183072];
  assign out_data[91583:91552] = in_data[183135:183104] - in_data[183167:183136];
  assign out_data[91615:91584] = in_data[183199:183168] - in_data[183231:183200];
  assign out_data[91647:91616] = in_data[183263:183232] - in_data[183295:183264];
  assign out_data[91679:91648] = in_data[183327:183296] - in_data[183359:183328];
  assign out_data[91711:91680] = in_data[183391:183360] - in_data[183423:183392];
  assign out_data[91743:91712] = in_data[183455:183424] - in_data[183487:183456];
  assign out_data[91775:91744] = in_data[183519:183488] - in_data[183551:183520];
  assign out_data[91807:91776] = in_data[183583:183552] - in_data[183615:183584];
  assign out_data[9183:9152] = in_data[18335:18304] - in_data[18367:18336];
  assign out_data[91839:91808] = in_data[183647:183616] - in_data[183679:183648];
  assign out_data[91871:91840] = in_data[183711:183680] - in_data[183743:183712];
  assign out_data[91903:91872] = in_data[183775:183744] - in_data[183807:183776];
  assign out_data[91935:91904] = in_data[183839:183808] - in_data[183871:183840];
  assign out_data[91967:91936] = in_data[183903:183872] - in_data[183935:183904];
  assign out_data[91999:91968] = in_data[183967:183936] - in_data[183999:183968];
  assign out_data[92031:92000] = in_data[184031:184000] - in_data[184063:184032];
  assign out_data[92063:92032] = in_data[184095:184064] - in_data[184127:184096];
  assign out_data[92095:92064] = in_data[184159:184128] - in_data[184191:184160];
  assign out_data[92127:92096] = in_data[184223:184192] - in_data[184255:184224];
  assign out_data[9215:9184] = in_data[18399:18368] - in_data[18431:18400];
  assign out_data[92159:92128] = in_data[184287:184256] - in_data[184319:184288];
  assign out_data[92191:92160] = in_data[184351:184320] - in_data[184383:184352];
  assign out_data[92223:92192] = in_data[184415:184384] - in_data[184447:184416];
  assign out_data[92255:92224] = in_data[184479:184448] - in_data[184511:184480];
  assign out_data[92287:92256] = in_data[184543:184512] - in_data[184575:184544];
  assign out_data[92319:92288] = in_data[184607:184576] - in_data[184639:184608];
  assign out_data[92351:92320] = in_data[184671:184640] - in_data[184703:184672];
  assign out_data[92383:92352] = in_data[184735:184704] - in_data[184767:184736];
  assign out_data[92415:92384] = in_data[184799:184768] - in_data[184831:184800];
  assign out_data[92447:92416] = in_data[184863:184832] - in_data[184895:184864];
  assign out_data[9247:9216] = in_data[18463:18432] - in_data[18495:18464];
  assign out_data[92479:92448] = in_data[184927:184896] - in_data[184959:184928];
  assign out_data[92511:92480] = in_data[184991:184960] - in_data[185023:184992];
  assign out_data[92543:92512] = in_data[185055:185024] - in_data[185087:185056];
  assign out_data[92575:92544] = in_data[185119:185088] - in_data[185151:185120];
  assign out_data[92607:92576] = in_data[185183:185152] - in_data[185215:185184];
  assign out_data[92639:92608] = in_data[185247:185216] - in_data[185279:185248];
  assign out_data[92671:92640] = in_data[185311:185280] - in_data[185343:185312];
  assign out_data[92703:92672] = in_data[185375:185344] - in_data[185407:185376];
  assign out_data[92735:92704] = in_data[185439:185408] - in_data[185471:185440];
  assign out_data[92767:92736] = in_data[185503:185472] - in_data[185535:185504];
  assign out_data[927:896] = in_data[1823:1792] - in_data[1855:1824];
  assign out_data[9279:9248] = in_data[18527:18496] - in_data[18559:18528];
  assign out_data[92799:92768] = in_data[185567:185536] - in_data[185599:185568];
  assign out_data[92831:92800] = in_data[185631:185600] - in_data[185663:185632];
  assign out_data[92863:92832] = in_data[185695:185664] - in_data[185727:185696];
  assign out_data[92895:92864] = in_data[185759:185728] - in_data[185791:185760];
  assign out_data[92927:92896] = in_data[185823:185792] - in_data[185855:185824];
  assign out_data[92959:92928] = in_data[185887:185856] - in_data[185919:185888];
  assign out_data[92991:92960] = in_data[185951:185920] - in_data[185983:185952];
  assign out_data[93023:92992] = in_data[186015:185984] - in_data[186047:186016];
  assign out_data[93055:93024] = in_data[186079:186048] - in_data[186111:186080];
  assign out_data[93087:93056] = in_data[186143:186112] - in_data[186175:186144];
  assign out_data[9311:9280] = in_data[18591:18560] - in_data[18623:18592];
  assign out_data[93119:93088] = in_data[186207:186176] - in_data[186239:186208];
  assign out_data[93151:93120] = in_data[186271:186240] - in_data[186303:186272];
  assign out_data[93183:93152] = in_data[186335:186304] - in_data[186367:186336];
  assign out_data[93215:93184] = in_data[186399:186368] - in_data[186431:186400];
  assign out_data[93247:93216] = in_data[186463:186432] - in_data[186495:186464];
  assign out_data[93279:93248] = in_data[186527:186496] - in_data[186559:186528];
  assign out_data[93311:93280] = in_data[186591:186560] - in_data[186623:186592];
  assign out_data[93343:93312] = in_data[186655:186624] - in_data[186687:186656];
  assign out_data[93375:93344] = in_data[186719:186688] - in_data[186751:186720];
  assign out_data[93407:93376] = in_data[186783:186752] - in_data[186815:186784];
  assign out_data[9343:9312] = in_data[18655:18624] - in_data[18687:18656];
  assign out_data[93439:93408] = in_data[186847:186816] - in_data[186879:186848];
  assign out_data[93471:93440] = in_data[186911:186880] - in_data[186943:186912];
  assign out_data[93503:93472] = in_data[186975:186944] - in_data[187007:186976];
  assign out_data[93535:93504] = in_data[187039:187008] - in_data[187071:187040];
  assign out_data[93567:93536] = in_data[187103:187072] - in_data[187135:187104];
  assign out_data[93599:93568] = in_data[187167:187136] - in_data[187199:187168];
  assign out_data[93631:93600] = in_data[187231:187200] - in_data[187263:187232];
  assign out_data[93663:93632] = in_data[187295:187264] - in_data[187327:187296];
  assign out_data[93695:93664] = in_data[187359:187328] - in_data[187391:187360];
  assign out_data[93727:93696] = in_data[187423:187392] - in_data[187455:187424];
  assign out_data[9375:9344] = in_data[18719:18688] - in_data[18751:18720];
  assign out_data[93759:93728] = in_data[187487:187456] - in_data[187519:187488];
  assign out_data[93791:93760] = in_data[187551:187520] - in_data[187583:187552];
  assign out_data[93823:93792] = in_data[187615:187584] - in_data[187647:187616];
  assign out_data[93855:93824] = in_data[187679:187648] - in_data[187711:187680];
  assign out_data[93887:93856] = in_data[187743:187712] - in_data[187775:187744];
  assign out_data[93919:93888] = in_data[187807:187776] - in_data[187839:187808];
  assign out_data[93951:93920] = in_data[187871:187840] - in_data[187903:187872];
  assign out_data[93983:93952] = in_data[187935:187904] - in_data[187967:187936];
  assign out_data[94015:93984] = in_data[187999:187968] - in_data[188031:188000];
  assign out_data[94047:94016] = in_data[188063:188032] - in_data[188095:188064];
  assign out_data[9407:9376] = in_data[18783:18752] - in_data[18815:18784];
  assign out_data[94079:94048] = in_data[188127:188096] - in_data[188159:188128];
  assign out_data[94111:94080] = in_data[188191:188160] - in_data[188223:188192];
  assign out_data[94143:94112] = in_data[188255:188224] - in_data[188287:188256];
  assign out_data[94175:94144] = in_data[188319:188288] - in_data[188351:188320];
  assign out_data[94207:94176] = in_data[188383:188352] - in_data[188415:188384];
  assign out_data[94239:94208] = in_data[188447:188416] - in_data[188479:188448];
  assign out_data[94271:94240] = in_data[188511:188480] - in_data[188543:188512];
  assign out_data[94303:94272] = in_data[188575:188544] - in_data[188607:188576];
  assign out_data[94335:94304] = in_data[188639:188608] - in_data[188671:188640];
  assign out_data[94367:94336] = in_data[188703:188672] - in_data[188735:188704];
  assign out_data[9439:9408] = in_data[18847:18816] - in_data[18879:18848];
  assign out_data[94399:94368] = in_data[188767:188736] - in_data[188799:188768];
  assign out_data[94431:94400] = in_data[188831:188800] - in_data[188863:188832];
  assign out_data[94463:94432] = in_data[188895:188864] - in_data[188927:188896];
  assign out_data[94495:94464] = in_data[188959:188928] - in_data[188991:188960];
  assign out_data[94527:94496] = in_data[189023:188992] - in_data[189055:189024];
  assign out_data[94559:94528] = in_data[189087:189056] - in_data[189119:189088];
  assign out_data[94591:94560] = in_data[189151:189120] - in_data[189183:189152];
  assign out_data[94623:94592] = in_data[189215:189184] - in_data[189247:189216];
  assign out_data[94655:94624] = in_data[189279:189248] - in_data[189311:189280];
  assign out_data[94687:94656] = in_data[189343:189312] - in_data[189375:189344];
  assign out_data[9471:9440] = in_data[18911:18880] - in_data[18943:18912];
  assign out_data[94719:94688] = in_data[189407:189376] - in_data[189439:189408];
  assign out_data[94751:94720] = in_data[189471:189440] - in_data[189503:189472];
  assign out_data[94783:94752] = in_data[189535:189504] - in_data[189567:189536];
  assign out_data[94815:94784] = in_data[189599:189568] - in_data[189631:189600];
  assign out_data[94847:94816] = in_data[189663:189632] - in_data[189695:189664];
  assign out_data[94879:94848] = in_data[189727:189696] - in_data[189759:189728];
  assign out_data[94911:94880] = in_data[189791:189760] - in_data[189823:189792];
  assign out_data[94943:94912] = in_data[189855:189824] - in_data[189887:189856];
  assign out_data[94975:94944] = in_data[189919:189888] - in_data[189951:189920];
  assign out_data[95007:94976] = in_data[189983:189952] - in_data[190015:189984];
  assign out_data[9503:9472] = in_data[18975:18944] - in_data[19007:18976];
  assign out_data[95039:95008] = in_data[190047:190016] - in_data[190079:190048];
  assign out_data[95071:95040] = in_data[190111:190080] - in_data[190143:190112];
  assign out_data[95103:95072] = in_data[190175:190144] - in_data[190207:190176];
  assign out_data[95135:95104] = in_data[190239:190208] - in_data[190271:190240];
  assign out_data[95167:95136] = in_data[190303:190272] - in_data[190335:190304];
  assign out_data[95199:95168] = in_data[190367:190336] - in_data[190399:190368];
  assign out_data[95231:95200] = in_data[190431:190400] - in_data[190463:190432];
  assign out_data[95263:95232] = in_data[190495:190464] - in_data[190527:190496];
  assign out_data[95295:95264] = in_data[190559:190528] - in_data[190591:190560];
  assign out_data[95327:95296] = in_data[190623:190592] - in_data[190655:190624];
  assign out_data[9535:9504] = in_data[19039:19008] - in_data[19071:19040];
  assign out_data[95359:95328] = in_data[190687:190656] - in_data[190719:190688];
  assign out_data[95391:95360] = in_data[190751:190720] - in_data[190783:190752];
  assign out_data[95423:95392] = in_data[190815:190784] - in_data[190847:190816];
  assign out_data[95455:95424] = in_data[190879:190848] - in_data[190911:190880];
  assign out_data[95487:95456] = in_data[190943:190912] - in_data[190975:190944];
  assign out_data[95519:95488] = in_data[191007:190976] - in_data[191039:191008];
  assign out_data[95551:95520] = in_data[191071:191040] - in_data[191103:191072];
  assign out_data[95583:95552] = in_data[191135:191104] - in_data[191167:191136];
  assign out_data[95615:95584] = in_data[191199:191168] - in_data[191231:191200];
  assign out_data[95647:95616] = in_data[191263:191232] - in_data[191295:191264];
  assign out_data[9567:9536] = in_data[19103:19072] - in_data[19135:19104];
  assign out_data[95679:95648] = in_data[191327:191296] - in_data[191359:191328];
  assign out_data[95711:95680] = in_data[191391:191360] - in_data[191423:191392];
  assign out_data[95743:95712] = in_data[191455:191424] - in_data[191487:191456];
  assign out_data[95775:95744] = in_data[191519:191488] - in_data[191551:191520];
  assign out_data[95807:95776] = in_data[191583:191552] - in_data[191615:191584];
  assign out_data[95839:95808] = in_data[191647:191616] - in_data[191679:191648];
  assign out_data[95871:95840] = in_data[191711:191680] - in_data[191743:191712];
  assign out_data[95903:95872] = in_data[191775:191744] - in_data[191807:191776];
  assign out_data[95935:95904] = in_data[191839:191808] - in_data[191871:191840];
  assign out_data[95967:95936] = in_data[191903:191872] - in_data[191935:191904];
  assign out_data[95:64] = in_data[159:128] - in_data[191:160];
  assign out_data[959:928] = in_data[1887:1856] - in_data[1919:1888];
  assign out_data[9599:9568] = in_data[19167:19136] - in_data[19199:19168];
  assign out_data[95999:95968] = in_data[191967:191936] - in_data[191999:191968];
  assign out_data[96031:96000] = in_data[192031:192000] - in_data[192063:192032];
  assign out_data[96063:96032] = in_data[192095:192064] - in_data[192127:192096];
  assign out_data[96095:96064] = in_data[192159:192128] - in_data[192191:192160];
  assign out_data[96127:96096] = in_data[192223:192192] - in_data[192255:192224];
  assign out_data[96159:96128] = in_data[192287:192256] - in_data[192319:192288];
  assign out_data[96191:96160] = in_data[192351:192320] - in_data[192383:192352];
  assign out_data[96223:96192] = in_data[192415:192384] - in_data[192447:192416];
  assign out_data[96255:96224] = in_data[192479:192448] - in_data[192511:192480];
  assign out_data[96287:96256] = in_data[192543:192512] - in_data[192575:192544];
  assign out_data[9631:9600] = in_data[19231:19200] - in_data[19263:19232];
  assign out_data[96319:96288] = in_data[192607:192576] - in_data[192639:192608];
  assign out_data[96351:96320] = in_data[192671:192640] - in_data[192703:192672];
  assign out_data[96383:96352] = in_data[192735:192704] - in_data[192767:192736];
  assign out_data[96415:96384] = in_data[192799:192768] - in_data[192831:192800];
  assign out_data[96447:96416] = in_data[192863:192832] - in_data[192895:192864];
  assign out_data[96479:96448] = in_data[192927:192896] - in_data[192959:192928];
  assign out_data[96511:96480] = in_data[192991:192960] - in_data[193023:192992];
  assign out_data[96543:96512] = in_data[193055:193024] - in_data[193087:193056];
  assign out_data[96575:96544] = in_data[193119:193088] - in_data[193151:193120];
  assign out_data[96607:96576] = in_data[193183:193152] - in_data[193215:193184];
  assign out_data[9663:9632] = in_data[19295:19264] - in_data[19327:19296];
  assign out_data[96639:96608] = in_data[193247:193216] - in_data[193279:193248];
  assign out_data[96671:96640] = in_data[193311:193280] - in_data[193343:193312];
  assign out_data[96703:96672] = in_data[193375:193344] - in_data[193407:193376];
  assign out_data[96735:96704] = in_data[193439:193408] - in_data[193471:193440];
  assign out_data[96767:96736] = in_data[193503:193472] - in_data[193535:193504];
  assign out_data[96799:96768] = in_data[193567:193536] - in_data[193599:193568];
  assign out_data[96831:96800] = in_data[193631:193600] - in_data[193663:193632];
  assign out_data[96863:96832] = in_data[193695:193664] - in_data[193727:193696];
  assign out_data[96895:96864] = in_data[193759:193728] - in_data[193791:193760];
  assign out_data[96927:96896] = in_data[193823:193792] - in_data[193855:193824];
  assign out_data[9695:9664] = in_data[19359:19328] - in_data[19391:19360];
  assign out_data[96959:96928] = in_data[193887:193856] - in_data[193919:193888];
  assign out_data[96991:96960] = in_data[193951:193920] - in_data[193983:193952];
  assign out_data[97023:96992] = in_data[194015:193984] - in_data[194047:194016];
  assign out_data[97055:97024] = in_data[194079:194048] - in_data[194111:194080];
  assign out_data[97087:97056] = in_data[194143:194112] - in_data[194175:194144];
  assign out_data[97119:97088] = in_data[194207:194176] - in_data[194239:194208];
  assign out_data[97151:97120] = in_data[194271:194240] - in_data[194303:194272];
  assign out_data[97183:97152] = in_data[194335:194304] - in_data[194367:194336];
  assign out_data[97215:97184] = in_data[194399:194368] - in_data[194431:194400];
  assign out_data[97247:97216] = in_data[194463:194432] - in_data[194495:194464];
  assign out_data[9727:9696] = in_data[19423:19392] - in_data[19455:19424];
  assign out_data[97279:97248] = in_data[194527:194496] - in_data[194559:194528];
  assign out_data[97311:97280] = in_data[194591:194560] - in_data[194623:194592];
  assign out_data[97343:97312] = in_data[194655:194624] - in_data[194687:194656];
  assign out_data[97375:97344] = in_data[194719:194688] - in_data[194751:194720];
  assign out_data[97407:97376] = in_data[194783:194752] - in_data[194815:194784];
  assign out_data[97439:97408] = in_data[194847:194816] - in_data[194879:194848];
  assign out_data[97471:97440] = in_data[194911:194880] - in_data[194943:194912];
  assign out_data[97503:97472] = in_data[194975:194944] - in_data[195007:194976];
  assign out_data[97535:97504] = in_data[195039:195008] - in_data[195071:195040];
  assign out_data[97567:97536] = in_data[195103:195072] - in_data[195135:195104];
  assign out_data[9759:9728] = in_data[19487:19456] - in_data[19519:19488];
  assign out_data[97599:97568] = in_data[195167:195136] - in_data[195199:195168];
  assign out_data[97631:97600] = in_data[195231:195200] - in_data[195263:195232];
  assign out_data[97663:97632] = in_data[195295:195264] - in_data[195327:195296];
  assign out_data[97695:97664] = in_data[195359:195328] - in_data[195391:195360];
  assign out_data[97727:97696] = in_data[195423:195392] - in_data[195455:195424];
  assign out_data[97759:97728] = in_data[195487:195456] - in_data[195519:195488];
  assign out_data[97791:97760] = in_data[195551:195520] - in_data[195583:195552];
  assign out_data[97823:97792] = in_data[195615:195584] - in_data[195647:195616];
  assign out_data[97855:97824] = in_data[195679:195648] - in_data[195711:195680];
  assign out_data[97887:97856] = in_data[195743:195712] - in_data[195775:195744];
  assign out_data[9791:9760] = in_data[19551:19520] - in_data[19583:19552];
  assign out_data[97919:97888] = in_data[195807:195776] - in_data[195839:195808];
  assign out_data[97951:97920] = in_data[195871:195840] - in_data[195903:195872];
  assign out_data[97983:97952] = in_data[195935:195904] - in_data[195967:195936];
  assign out_data[98015:97984] = in_data[195999:195968] - in_data[196031:196000];
  assign out_data[98047:98016] = in_data[196063:196032] - in_data[196095:196064];
  assign out_data[98079:98048] = in_data[196127:196096] - in_data[196159:196128];
  assign out_data[98111:98080] = in_data[196191:196160] - in_data[196223:196192];
  assign out_data[98143:98112] = in_data[196255:196224] - in_data[196287:196256];
  assign out_data[98175:98144] = in_data[196319:196288] - in_data[196351:196320];
  assign out_data[98207:98176] = in_data[196383:196352] - in_data[196415:196384];
  assign out_data[9823:9792] = in_data[19615:19584] - in_data[19647:19616];
  assign out_data[98239:98208] = in_data[196447:196416] - in_data[196479:196448];
  assign out_data[98271:98240] = in_data[196511:196480] - in_data[196543:196512];
  assign out_data[98303:98272] = in_data[196575:196544] - in_data[196607:196576];
  assign out_data[98335:98304] = in_data[196639:196608] - in_data[196671:196640];
  assign out_data[98367:98336] = in_data[196703:196672] - in_data[196735:196704];
  assign out_data[98399:98368] = in_data[196767:196736] - in_data[196799:196768];
  assign out_data[98431:98400] = in_data[196831:196800] - in_data[196863:196832];
  assign out_data[98463:98432] = in_data[196895:196864] - in_data[196927:196896];
  assign out_data[98495:98464] = in_data[196959:196928] - in_data[196991:196960];
  assign out_data[98527:98496] = in_data[197023:196992] - in_data[197055:197024];
  assign out_data[9855:9824] = in_data[19679:19648] - in_data[19711:19680];
  assign out_data[98559:98528] = in_data[197087:197056] - in_data[197119:197088];
  assign out_data[98591:98560] = in_data[197151:197120] - in_data[197183:197152];
  assign out_data[98623:98592] = in_data[197215:197184] - in_data[197247:197216];
  assign out_data[98655:98624] = in_data[197279:197248] - in_data[197311:197280];
  assign out_data[98687:98656] = in_data[197343:197312] - in_data[197375:197344];
  assign out_data[98719:98688] = in_data[197407:197376] - in_data[197439:197408];
  assign out_data[98751:98720] = in_data[197471:197440] - in_data[197503:197472];
  assign out_data[98783:98752] = in_data[197535:197504] - in_data[197567:197536];
  assign out_data[98815:98784] = in_data[197599:197568] - in_data[197631:197600];
  assign out_data[98847:98816] = in_data[197663:197632] - in_data[197695:197664];
  assign out_data[9887:9856] = in_data[19743:19712] - in_data[19775:19744];
  assign out_data[98879:98848] = in_data[197727:197696] - in_data[197759:197728];
  assign out_data[98911:98880] = in_data[197791:197760] - in_data[197823:197792];
  assign out_data[98943:98912] = in_data[197855:197824] - in_data[197887:197856];
  assign out_data[98975:98944] = in_data[197919:197888] - in_data[197951:197920];
  assign out_data[99007:98976] = in_data[197983:197952] - in_data[198015:197984];
  assign out_data[99039:99008] = in_data[198047:198016] - in_data[198079:198048];
  assign out_data[99071:99040] = in_data[198111:198080] - in_data[198143:198112];
  assign out_data[99103:99072] = in_data[198175:198144] - in_data[198207:198176];
  assign out_data[99135:99104] = in_data[198239:198208] - in_data[198271:198240];
  assign out_data[99167:99136] = in_data[198303:198272] - in_data[198335:198304];
  assign out_data[991:960] = in_data[1951:1920] - in_data[1983:1952];
  assign out_data[9919:9888] = in_data[19807:19776] - in_data[19839:19808];
  assign out_data[99199:99168] = in_data[198367:198336] - in_data[198399:198368];
  assign out_data[99231:99200] = in_data[198431:198400] - in_data[198463:198432];
  assign out_data[99263:99232] = in_data[198495:198464] - in_data[198527:198496];
  assign out_data[99295:99264] = in_data[198559:198528] - in_data[198591:198560];
  assign out_data[99327:99296] = in_data[198623:198592] - in_data[198655:198624];
  assign out_data[99359:99328] = in_data[198687:198656] - in_data[198719:198688];
  assign out_data[99391:99360] = in_data[198751:198720] - in_data[198783:198752];
  assign out_data[99423:99392] = in_data[198815:198784] - in_data[198847:198816];
  assign out_data[99455:99424] = in_data[198879:198848] - in_data[198911:198880];
  assign out_data[99487:99456] = in_data[198943:198912] - in_data[198975:198944];
  assign out_data[9951:9920] = in_data[19871:19840] - in_data[19903:19872];
  assign out_data[99519:99488] = in_data[199007:198976] - in_data[199039:199008];
  assign out_data[99551:99520] = in_data[199071:199040] - in_data[199103:199072];
  assign out_data[99583:99552] = in_data[199135:199104] - in_data[199167:199136];
  assign out_data[99615:99584] = in_data[199199:199168] - in_data[199231:199200];
  assign out_data[99647:99616] = in_data[199263:199232] - in_data[199295:199264];
  assign out_data[99679:99648] = in_data[199327:199296] - in_data[199359:199328];
  assign out_data[99711:99680] = in_data[199391:199360] - in_data[199423:199392];
  assign out_data[99743:99712] = in_data[199455:199424] - in_data[199487:199456];
  assign out_data[99775:99744] = in_data[199519:199488] - in_data[199551:199520];
  assign out_data[99807:99776] = in_data[199583:199552] - in_data[199615:199584];
  assign out_data[9983:9952] = in_data[19935:19904] - in_data[19967:19936];
  assign out_data[99839:99808] = in_data[199647:199616] - in_data[199679:199648];
  assign out_data[99871:99840] = in_data[199711:199680] - in_data[199743:199712];
  assign out_data[99903:99872] = in_data[199775:199744] - in_data[199807:199776];
  assign out_data[99935:99904] = in_data[199839:199808] - in_data[199871:199840];
  assign out_data[99967:99936] = in_data[199903:199872] - in_data[199935:199904];
  assign out_data[99999:99968] = in_data[199967:199936] - in_data[199999:199968];
  assign out_data[100031:100000] = in_data[200031:200000] - in_data[200063:200032];
  assign out_data[100063:100032] = in_data[200095:200064] - in_data[200127:200096];
  assign out_data[100095:100064] = in_data[200159:200128] - in_data[200191:200160];
  assign out_data[100127:100096] = in_data[200223:200192] - in_data[200255:200224];
  assign out_data[10015:9984] = in_data[19999:19968] - in_data[20031:20000];
  assign out_data[100159:100128] = in_data[200287:200256] - in_data[200319:200288];
  assign out_data[100191:100160] = in_data[200351:200320] - in_data[200383:200352];
  assign out_data[100223:100192] = in_data[200415:200384] - in_data[200447:200416];
  assign out_data[100255:100224] = in_data[200479:200448] - in_data[200511:200480];
  assign out_data[100287:100256] = in_data[200543:200512] - in_data[200575:200544];
  assign out_data[100319:100288] = in_data[200607:200576] - in_data[200639:200608];
  assign out_data[100351:100320] = in_data[200671:200640] - in_data[200703:200672];
  assign out_data[100383:100352] = in_data[200735:200704] - in_data[200767:200736];
  assign out_data[100415:100384] = in_data[200799:200768] - in_data[200831:200800];
  assign out_data[100447:100416] = in_data[200863:200832] - in_data[200895:200864];
  assign out_data[10047:10016] = in_data[20063:20032] - in_data[20095:20064];
  assign out_data[100479:100448] = in_data[200927:200896] - in_data[200959:200928];
  assign out_data[100511:100480] = in_data[200991:200960] - in_data[201023:200992];
  assign out_data[100543:100512] = in_data[201055:201024] - in_data[201087:201056];
  assign out_data[100575:100544] = in_data[201119:201088] - in_data[201151:201120];
  assign out_data[100607:100576] = in_data[201183:201152] - in_data[201215:201184];
  assign out_data[100639:100608] = in_data[201247:201216] - in_data[201279:201248];
  assign out_data[100671:100640] = in_data[201311:201280] - in_data[201343:201312];
  assign out_data[100703:100672] = in_data[201375:201344] - in_data[201407:201376];
  assign out_data[100735:100704] = in_data[201439:201408] - in_data[201471:201440];
  assign out_data[100767:100736] = in_data[201503:201472] - in_data[201535:201504];
  assign out_data[10079:10048] = in_data[20127:20096] - in_data[20159:20128];
  assign out_data[100799:100768] = in_data[201567:201536] - in_data[201599:201568];
  assign out_data[100831:100800] = in_data[201631:201600] - in_data[201663:201632];
  assign out_data[100863:100832] = in_data[201695:201664] - in_data[201727:201696];
  assign out_data[100895:100864] = in_data[201759:201728] - in_data[201791:201760];
  assign out_data[100927:100896] = in_data[201823:201792] - in_data[201855:201824];
  assign out_data[100959:100928] = in_data[201887:201856] - in_data[201919:201888];
  assign out_data[100991:100960] = in_data[201951:201920] - in_data[201983:201952];
  assign out_data[101023:100992] = in_data[202015:201984] - in_data[202047:202016];
  assign out_data[101055:101024] = in_data[202079:202048] - in_data[202111:202080];
  assign out_data[101087:101056] = in_data[202143:202112] - in_data[202175:202144];
  assign out_data[10111:10080] = in_data[20191:20160] - in_data[20223:20192];
  assign out_data[101119:101088] = in_data[202207:202176] - in_data[202239:202208];
  assign out_data[101151:101120] = in_data[202271:202240] - in_data[202303:202272];
  assign out_data[101183:101152] = in_data[202335:202304] - in_data[202367:202336];
  assign out_data[101215:101184] = in_data[202399:202368] - in_data[202431:202400];
  assign out_data[101247:101216] = in_data[202463:202432] - in_data[202495:202464];
  assign out_data[101279:101248] = in_data[202527:202496] - in_data[202559:202528];
  assign out_data[101311:101280] = in_data[202591:202560] - in_data[202623:202592];
  assign out_data[101343:101312] = in_data[202655:202624] - in_data[202687:202656];
  assign out_data[101375:101344] = in_data[202719:202688] - in_data[202751:202720];
  assign out_data[101407:101376] = in_data[202783:202752] - in_data[202815:202784];
  assign out_data[10143:10112] = in_data[20255:20224] - in_data[20287:20256];
  assign out_data[101439:101408] = in_data[202847:202816] - in_data[202879:202848];
  assign out_data[101471:101440] = in_data[202911:202880] - in_data[202943:202912];
  assign out_data[101503:101472] = in_data[202975:202944] - in_data[203007:202976];
  assign out_data[101535:101504] = in_data[203039:203008] - in_data[203071:203040];
  assign out_data[101567:101536] = in_data[203103:203072] - in_data[203135:203104];
  assign out_data[101599:101568] = in_data[203167:203136] - in_data[203199:203168];
  assign out_data[101631:101600] = in_data[203231:203200] - in_data[203263:203232];
  assign out_data[101663:101632] = in_data[203295:203264] - in_data[203327:203296];
  assign out_data[101695:101664] = in_data[203359:203328] - in_data[203391:203360];
  assign out_data[101727:101696] = in_data[203423:203392] - in_data[203455:203424];
  assign out_data[10175:10144] = in_data[20319:20288] - in_data[20351:20320];
  assign out_data[101759:101728] = in_data[203487:203456] - in_data[203519:203488];
  assign out_data[101791:101760] = in_data[203551:203520] - in_data[203583:203552];
  assign out_data[101823:101792] = in_data[203615:203584] - in_data[203647:203616];
  assign out_data[101855:101824] = in_data[203679:203648] - in_data[203711:203680];
  assign out_data[101887:101856] = in_data[203743:203712] - in_data[203775:203744];
  assign out_data[101919:101888] = in_data[203807:203776] - in_data[203839:203808];
  assign out_data[101951:101920] = in_data[203871:203840] - in_data[203903:203872];
  assign out_data[101983:101952] = in_data[203935:203904] - in_data[203967:203936];
  assign out_data[102015:101984] = in_data[203999:203968] - in_data[204031:204000];
  assign out_data[102047:102016] = in_data[204063:204032] - in_data[204095:204064];
  assign out_data[10207:10176] = in_data[20383:20352] - in_data[20415:20384];
  assign out_data[102079:102048] = in_data[204127:204096] - in_data[204159:204128];
  assign out_data[102111:102080] = in_data[204191:204160] - in_data[204223:204192];
  assign out_data[102143:102112] = in_data[204255:204224] - in_data[204287:204256];
  assign out_data[102175:102144] = in_data[204319:204288] - in_data[204351:204320];
  assign out_data[102207:102176] = in_data[204383:204352] - in_data[204415:204384];
  assign out_data[102239:102208] = in_data[204447:204416] - in_data[204479:204448];
  assign out_data[102271:102240] = in_data[204511:204480] - in_data[204543:204512];
  assign out_data[102303:102272] = in_data[204575:204544] - in_data[204607:204576];
  assign out_data[102335:102304] = in_data[204639:204608] - in_data[204671:204640];
  assign out_data[102367:102336] = in_data[204703:204672] - in_data[204735:204704];
  assign out_data[1023:992] = in_data[2015:1984] - in_data[2047:2016];
  assign out_data[10239:10208] = in_data[20447:20416] - in_data[20479:20448];
  assign out_data[102399:102368] = in_data[204767:204736] - in_data[204799:204768];
  assign out_data[102431:102400] = in_data[204831:204800] - in_data[204863:204832];
  assign out_data[102463:102432] = in_data[204895:204864] - in_data[204927:204896];
  assign out_data[102495:102464] = in_data[204959:204928] - in_data[204991:204960];
  assign out_data[102527:102496] = in_data[205023:204992] - in_data[205055:205024];
  assign out_data[102559:102528] = in_data[205087:205056] - in_data[205119:205088];
  assign out_data[102591:102560] = in_data[205151:205120] - in_data[205183:205152];
  assign out_data[102623:102592] = in_data[205215:205184] - in_data[205247:205216];
  assign out_data[102655:102624] = in_data[205279:205248] - in_data[205311:205280];
  assign out_data[102687:102656] = in_data[205343:205312] - in_data[205375:205344];
  assign out_data[10271:10240] = in_data[20511:20480] - in_data[20543:20512];
  assign out_data[102719:102688] = in_data[205407:205376] - in_data[205439:205408];
  assign out_data[102751:102720] = in_data[205471:205440] - in_data[205503:205472];
  assign out_data[102783:102752] = in_data[205535:205504] - in_data[205567:205536];
  assign out_data[102815:102784] = in_data[205599:205568] - in_data[205631:205600];
  assign out_data[102847:102816] = in_data[205663:205632] - in_data[205695:205664];
  assign out_data[102879:102848] = in_data[205727:205696] - in_data[205759:205728];
  assign out_data[102911:102880] = in_data[205791:205760] - in_data[205823:205792];
  assign out_data[102943:102912] = in_data[205855:205824] - in_data[205887:205856];
  assign out_data[102975:102944] = in_data[205919:205888] - in_data[205951:205920];
  assign out_data[103007:102976] = in_data[205983:205952] - in_data[206015:205984];
  assign out_data[10303:10272] = in_data[20575:20544] - in_data[20607:20576];
  assign out_data[103039:103008] = in_data[206047:206016] - in_data[206079:206048];
  assign out_data[103071:103040] = in_data[206111:206080] - in_data[206143:206112];
  assign out_data[103103:103072] = in_data[206175:206144] - in_data[206207:206176];
  assign out_data[103135:103104] = in_data[206239:206208] - in_data[206271:206240];
  assign out_data[103167:103136] = in_data[206303:206272] - in_data[206335:206304];
  assign out_data[103199:103168] = in_data[206367:206336] - in_data[206399:206368];
  assign out_data[103231:103200] = in_data[206431:206400] - in_data[206463:206432];
  assign out_data[103263:103232] = in_data[206495:206464] - in_data[206527:206496];
  assign out_data[103295:103264] = in_data[206559:206528] - in_data[206591:206560];
  assign out_data[103327:103296] = in_data[206623:206592] - in_data[206655:206624];
  assign out_data[10335:10304] = in_data[20639:20608] - in_data[20671:20640];
  assign out_data[103359:103328] = in_data[206687:206656] - in_data[206719:206688];
  assign out_data[103391:103360] = in_data[206751:206720] - in_data[206783:206752];
  assign out_data[103423:103392] = in_data[206815:206784] - in_data[206847:206816];
  assign out_data[103455:103424] = in_data[206879:206848] - in_data[206911:206880];
  assign out_data[103487:103456] = in_data[206943:206912] - in_data[206975:206944];
  assign out_data[103519:103488] = in_data[207007:206976] - in_data[207039:207008];
  assign out_data[103551:103520] = in_data[207071:207040] - in_data[207103:207072];
  assign out_data[103583:103552] = in_data[207135:207104] - in_data[207167:207136];
  assign out_data[103615:103584] = in_data[207199:207168] - in_data[207231:207200];
  assign out_data[103647:103616] = in_data[207263:207232] - in_data[207295:207264];
  assign out_data[10367:10336] = in_data[20703:20672] - in_data[20735:20704];
  assign out_data[103679:103648] = in_data[207327:207296] - in_data[207359:207328];
  assign out_data[103711:103680] = in_data[207391:207360] - in_data[207423:207392];
  assign out_data[103743:103712] = in_data[207455:207424] - in_data[207487:207456];
  assign out_data[103775:103744] = in_data[207519:207488] - in_data[207551:207520];
  assign out_data[103807:103776] = in_data[207583:207552] - in_data[207615:207584];
  assign out_data[103839:103808] = in_data[207647:207616] - in_data[207679:207648];
  assign out_data[103871:103840] = in_data[207711:207680] - in_data[207743:207712];
  assign out_data[103903:103872] = in_data[207775:207744] - in_data[207807:207776];
  assign out_data[103935:103904] = in_data[207839:207808] - in_data[207871:207840];
  assign out_data[103967:103936] = in_data[207903:207872] - in_data[207935:207904];
  assign out_data[10399:10368] = in_data[20767:20736] - in_data[20799:20768];
  assign out_data[103999:103968] = in_data[207967:207936] - in_data[207999:207968];
  assign out_data[104031:104000] = in_data[208031:208000] - in_data[208063:208032];
  assign out_data[104063:104032] = in_data[208095:208064] - in_data[208127:208096];
  assign out_data[104095:104064] = in_data[208159:208128] - in_data[208191:208160];
  assign out_data[104127:104096] = in_data[208223:208192] - in_data[208255:208224];
  assign out_data[104159:104128] = in_data[208287:208256] - in_data[208319:208288];
  assign out_data[104191:104160] = in_data[208351:208320] - in_data[208383:208352];
  assign out_data[104223:104192] = in_data[208415:208384] - in_data[208447:208416];
  assign out_data[104255:104224] = in_data[208479:208448] - in_data[208511:208480];
  assign out_data[104287:104256] = in_data[208543:208512] - in_data[208575:208544];
  assign out_data[10431:10400] = in_data[20831:20800] - in_data[20863:20832];
  assign out_data[104319:104288] = in_data[208607:208576] - in_data[208639:208608];
  assign out_data[104351:104320] = in_data[208671:208640] - in_data[208703:208672];
  assign out_data[104383:104352] = in_data[208735:208704] - in_data[208767:208736];
  assign out_data[104415:104384] = in_data[208799:208768] - in_data[208831:208800];
  assign out_data[104447:104416] = in_data[208863:208832] - in_data[208895:208864];
  assign out_data[104479:104448] = in_data[208927:208896] - in_data[208959:208928];
  assign out_data[104511:104480] = in_data[208991:208960] - in_data[209023:208992];
  assign out_data[104543:104512] = in_data[209055:209024] - in_data[209087:209056];
  assign out_data[104575:104544] = in_data[209119:209088] - in_data[209151:209120];
  assign out_data[104607:104576] = in_data[209183:209152] - in_data[209215:209184];
  assign out_data[10463:10432] = in_data[20895:20864] - in_data[20927:20896];
  assign out_data[104639:104608] = in_data[209247:209216] - in_data[209279:209248];
  assign out_data[104671:104640] = in_data[209311:209280] - in_data[209343:209312];
  assign out_data[104703:104672] = in_data[209375:209344] - in_data[209407:209376];
  assign out_data[104735:104704] = in_data[209439:209408] - in_data[209471:209440];
  assign out_data[104767:104736] = in_data[209503:209472] - in_data[209535:209504];
  assign out_data[104799:104768] = in_data[209567:209536] - in_data[209599:209568];
  assign out_data[104831:104800] = in_data[209631:209600] - in_data[209663:209632];
  assign out_data[104863:104832] = in_data[209695:209664] - in_data[209727:209696];
  assign out_data[104895:104864] = in_data[209759:209728] - in_data[209791:209760];
  assign out_data[104927:104896] = in_data[209823:209792] - in_data[209855:209824];
  assign out_data[10495:10464] = in_data[20959:20928] - in_data[20991:20960];
  assign out_data[104959:104928] = in_data[209887:209856] - in_data[209919:209888];
  assign out_data[104991:104960] = in_data[209951:209920] - in_data[209983:209952];
  assign out_data[105023:104992] = in_data[210015:209984] - in_data[210047:210016];
  assign out_data[105055:105024] = in_data[210079:210048] - in_data[210111:210080];
  assign out_data[105087:105056] = in_data[210143:210112] - in_data[210175:210144];
  assign out_data[105119:105088] = in_data[210207:210176] - in_data[210239:210208];
  assign out_data[105151:105120] = in_data[210271:210240] - in_data[210303:210272];
  assign out_data[105183:105152] = in_data[210335:210304] - in_data[210367:210336];
  assign out_data[105215:105184] = in_data[210399:210368] - in_data[210431:210400];
  assign out_data[105247:105216] = in_data[210463:210432] - in_data[210495:210464];
  assign out_data[10527:10496] = in_data[21023:20992] - in_data[21055:21024];
  assign out_data[105279:105248] = in_data[210527:210496] - in_data[210559:210528];
  assign out_data[105311:105280] = in_data[210591:210560] - in_data[210623:210592];
  assign out_data[105343:105312] = in_data[210655:210624] - in_data[210687:210656];
  assign out_data[105375:105344] = in_data[210719:210688] - in_data[210751:210720];
  assign out_data[105407:105376] = in_data[210783:210752] - in_data[210815:210784];
  assign out_data[105439:105408] = in_data[210847:210816] - in_data[210879:210848];
  assign out_data[105471:105440] = in_data[210911:210880] - in_data[210943:210912];
  assign out_data[105503:105472] = in_data[210975:210944] - in_data[211007:210976];
  assign out_data[105535:105504] = in_data[211039:211008] - in_data[211071:211040];
  assign out_data[105567:105536] = in_data[211103:211072] - in_data[211135:211104];
  assign out_data[1055:1024] = in_data[2079:2048] - in_data[2111:2080];
  assign out_data[10559:10528] = in_data[21087:21056] - in_data[21119:21088];
  assign out_data[105599:105568] = in_data[211167:211136] - in_data[211199:211168];
  assign out_data[105631:105600] = in_data[211231:211200] - in_data[211263:211232];
  assign out_data[105663:105632] = in_data[211295:211264] - in_data[211327:211296];
  assign out_data[105695:105664] = in_data[211359:211328] - in_data[211391:211360];
  assign out_data[105727:105696] = in_data[211423:211392] - in_data[211455:211424];
  assign out_data[105759:105728] = in_data[211487:211456] - in_data[211519:211488];
  assign out_data[105791:105760] = in_data[211551:211520] - in_data[211583:211552];
  assign out_data[105823:105792] = in_data[211615:211584] - in_data[211647:211616];
  assign out_data[105855:105824] = in_data[211679:211648] - in_data[211711:211680];
  assign out_data[105887:105856] = in_data[211743:211712] - in_data[211775:211744];
  assign out_data[10591:10560] = in_data[21151:21120] - in_data[21183:21152];
  assign out_data[105919:105888] = in_data[211807:211776] - in_data[211839:211808];
  assign out_data[105951:105920] = in_data[211871:211840] - in_data[211903:211872];
  assign out_data[105983:105952] = in_data[211935:211904] - in_data[211967:211936];
  assign out_data[106015:105984] = in_data[211999:211968] - in_data[212031:212000];
  assign out_data[106047:106016] = in_data[212063:212032] - in_data[212095:212064];
  assign out_data[106079:106048] = in_data[212127:212096] - in_data[212159:212128];
  assign out_data[106111:106080] = in_data[212191:212160] - in_data[212223:212192];
  assign out_data[106143:106112] = in_data[212255:212224] - in_data[212287:212256];
  assign out_data[106175:106144] = in_data[212319:212288] - in_data[212351:212320];
  assign out_data[106207:106176] = in_data[212383:212352] - in_data[212415:212384];
  assign out_data[10623:10592] = in_data[21215:21184] - in_data[21247:21216];
  assign out_data[106239:106208] = in_data[212447:212416] - in_data[212479:212448];
  assign out_data[106271:106240] = in_data[212511:212480] - in_data[212543:212512];
  assign out_data[106303:106272] = in_data[212575:212544] - in_data[212607:212576];
  assign out_data[106335:106304] = in_data[212639:212608] - in_data[212671:212640];
  assign out_data[106367:106336] = in_data[212703:212672] - in_data[212735:212704];
  assign out_data[106399:106368] = in_data[212767:212736] - in_data[212799:212768];
  assign out_data[106431:106400] = in_data[212831:212800] - in_data[212863:212832];
  assign out_data[106463:106432] = in_data[212895:212864] - in_data[212927:212896];
  assign out_data[106495:106464] = in_data[212959:212928] - in_data[212991:212960];
  assign out_data[106527:106496] = in_data[213023:212992] - in_data[213055:213024];
  assign out_data[10655:10624] = in_data[21279:21248] - in_data[21311:21280];
  assign out_data[106559:106528] = in_data[213087:213056] - in_data[213119:213088];
  assign out_data[106591:106560] = in_data[213151:213120] - in_data[213183:213152];
  assign out_data[106623:106592] = in_data[213215:213184] - in_data[213247:213216];
  assign out_data[106655:106624] = in_data[213279:213248] - in_data[213311:213280];
  assign out_data[106687:106656] = in_data[213343:213312] - in_data[213375:213344];
  assign out_data[106719:106688] = in_data[213407:213376] - in_data[213439:213408];
  assign out_data[106751:106720] = in_data[213471:213440] - in_data[213503:213472];
  assign out_data[106783:106752] = in_data[213535:213504] - in_data[213567:213536];
  assign out_data[106815:106784] = in_data[213599:213568] - in_data[213631:213600];
  assign out_data[106847:106816] = in_data[213663:213632] - in_data[213695:213664];
  assign out_data[10687:10656] = in_data[21343:21312] - in_data[21375:21344];
  assign out_data[106879:106848] = in_data[213727:213696] - in_data[213759:213728];
  assign out_data[106911:106880] = in_data[213791:213760] - in_data[213823:213792];
  assign out_data[106943:106912] = in_data[213855:213824] - in_data[213887:213856];
  assign out_data[106975:106944] = in_data[213919:213888] - in_data[213951:213920];
  assign out_data[107007:106976] = in_data[213983:213952] - in_data[214015:213984];
  assign out_data[107039:107008] = in_data[214047:214016] - in_data[214079:214048];
  assign out_data[107071:107040] = in_data[214111:214080] - in_data[214143:214112];
  assign out_data[107103:107072] = in_data[214175:214144] - in_data[214207:214176];
  assign out_data[107135:107104] = in_data[214239:214208] - in_data[214271:214240];
  assign out_data[107167:107136] = in_data[214303:214272] - in_data[214335:214304];
  assign out_data[10719:10688] = in_data[21407:21376] - in_data[21439:21408];
  assign out_data[107199:107168] = in_data[214367:214336] - in_data[214399:214368];
  assign out_data[107231:107200] = in_data[214431:214400] - in_data[214463:214432];
  assign out_data[107263:107232] = in_data[214495:214464] - in_data[214527:214496];
  assign out_data[107295:107264] = in_data[214559:214528] - in_data[214591:214560];
  assign out_data[107327:107296] = in_data[214623:214592] - in_data[214655:214624];
  assign out_data[107359:107328] = in_data[214687:214656] - in_data[214719:214688];
  assign out_data[107391:107360] = in_data[214751:214720] - in_data[214783:214752];
  assign out_data[107423:107392] = in_data[214815:214784] - in_data[214847:214816];
  assign out_data[107455:107424] = in_data[214879:214848] - in_data[214911:214880];
  assign out_data[107487:107456] = in_data[214943:214912] - in_data[214975:214944];
  assign out_data[10751:10720] = in_data[21471:21440] - in_data[21503:21472];
  assign out_data[107519:107488] = in_data[215007:214976] - in_data[215039:215008];
  assign out_data[107551:107520] = in_data[215071:215040] - in_data[215103:215072];
  assign out_data[107583:107552] = in_data[215135:215104] - in_data[215167:215136];
  assign out_data[107615:107584] = in_data[215199:215168] - in_data[215231:215200];
  assign out_data[107647:107616] = in_data[215263:215232] - in_data[215295:215264];
  assign out_data[107679:107648] = in_data[215327:215296] - in_data[215359:215328];
  assign out_data[107711:107680] = in_data[215391:215360] - in_data[215423:215392];
  assign out_data[107743:107712] = in_data[215455:215424] - in_data[215487:215456];
  assign out_data[107775:107744] = in_data[215519:215488] - in_data[215551:215520];
  assign out_data[107807:107776] = in_data[215583:215552] - in_data[215615:215584];
  assign out_data[10783:10752] = in_data[21535:21504] - in_data[21567:21536];
  assign out_data[107839:107808] = in_data[215647:215616] - in_data[215679:215648];
  assign out_data[107871:107840] = in_data[215711:215680] - in_data[215743:215712];
  assign out_data[107903:107872] = in_data[215775:215744] - in_data[215807:215776];
  assign out_data[107935:107904] = in_data[215839:215808] - in_data[215871:215840];
  assign out_data[107967:107936] = in_data[215903:215872] - in_data[215935:215904];
  assign out_data[107999:107968] = in_data[215967:215936] - in_data[215999:215968];
  assign out_data[108031:108000] = in_data[216031:216000] - in_data[216063:216032];
  assign out_data[108063:108032] = in_data[216095:216064] - in_data[216127:216096];
  assign out_data[108095:108064] = in_data[216159:216128] - in_data[216191:216160];
  assign out_data[108127:108096] = in_data[216223:216192] - in_data[216255:216224];
  assign out_data[10815:10784] = in_data[21599:21568] - in_data[21631:21600];
  assign out_data[108159:108128] = in_data[216287:216256] - in_data[216319:216288];
  assign out_data[108191:108160] = in_data[216351:216320] - in_data[216383:216352];
  assign out_data[108223:108192] = in_data[216415:216384] - in_data[216447:216416];
  assign out_data[108255:108224] = in_data[216479:216448] - in_data[216511:216480];
  assign out_data[108287:108256] = in_data[216543:216512] - in_data[216575:216544];
  assign out_data[108319:108288] = in_data[216607:216576] - in_data[216639:216608];
  assign out_data[108351:108320] = in_data[216671:216640] - in_data[216703:216672];
  assign out_data[108383:108352] = in_data[216735:216704] - in_data[216767:216736];
  assign out_data[108415:108384] = in_data[216799:216768] - in_data[216831:216800];
  assign out_data[108447:108416] = in_data[216863:216832] - in_data[216895:216864];
  assign out_data[10847:10816] = in_data[21663:21632] - in_data[21695:21664];
  assign out_data[108479:108448] = in_data[216927:216896] - in_data[216959:216928];
  assign out_data[108511:108480] = in_data[216991:216960] - in_data[217023:216992];
  assign out_data[108543:108512] = in_data[217055:217024] - in_data[217087:217056];
  assign out_data[108575:108544] = in_data[217119:217088] - in_data[217151:217120];
  assign out_data[108607:108576] = in_data[217183:217152] - in_data[217215:217184];
  assign out_data[108639:108608] = in_data[217247:217216] - in_data[217279:217248];
  assign out_data[108671:108640] = in_data[217311:217280] - in_data[217343:217312];
  assign out_data[108703:108672] = in_data[217375:217344] - in_data[217407:217376];
  assign out_data[108735:108704] = in_data[217439:217408] - in_data[217471:217440];
  assign out_data[108767:108736] = in_data[217503:217472] - in_data[217535:217504];
  assign out_data[1087:1056] = in_data[2143:2112] - in_data[2175:2144];
  assign out_data[10879:10848] = in_data[21727:21696] - in_data[21759:21728];
  assign out_data[108799:108768] = in_data[217567:217536] - in_data[217599:217568];
  assign out_data[108831:108800] = in_data[217631:217600] - in_data[217663:217632];
  assign out_data[108863:108832] = in_data[217695:217664] - in_data[217727:217696];
  assign out_data[108895:108864] = in_data[217759:217728] - in_data[217791:217760];
  assign out_data[108927:108896] = in_data[217823:217792] - in_data[217855:217824];
  assign out_data[108959:108928] = in_data[217887:217856] - in_data[217919:217888];
  assign out_data[108991:108960] = in_data[217951:217920] - in_data[217983:217952];
  assign out_data[109023:108992] = in_data[218015:217984] - in_data[218047:218016];
  assign out_data[109055:109024] = in_data[218079:218048] - in_data[218111:218080];
  assign out_data[109087:109056] = in_data[218143:218112] - in_data[218175:218144];
  assign out_data[10911:10880] = in_data[21791:21760] - in_data[21823:21792];
  assign out_data[109119:109088] = in_data[218207:218176] - in_data[218239:218208];
  assign out_data[109151:109120] = in_data[218271:218240] - in_data[218303:218272];
  assign out_data[109183:109152] = in_data[218335:218304] - in_data[218367:218336];
  assign out_data[109215:109184] = in_data[218399:218368] - in_data[218431:218400];
  assign out_data[109247:109216] = in_data[218463:218432] - in_data[218495:218464];
  assign out_data[109279:109248] = in_data[218527:218496] - in_data[218559:218528];
  assign out_data[109311:109280] = in_data[218591:218560] - in_data[218623:218592];
  assign out_data[109343:109312] = in_data[218655:218624] - in_data[218687:218656];
  assign out_data[109375:109344] = in_data[218719:218688] - in_data[218751:218720];
  assign out_data[109407:109376] = in_data[218783:218752] - in_data[218815:218784];
  assign out_data[10943:10912] = in_data[21855:21824] - in_data[21887:21856];
  assign out_data[109439:109408] = in_data[218847:218816] - in_data[218879:218848];
  assign out_data[109471:109440] = in_data[218911:218880] - in_data[218943:218912];
  assign out_data[109503:109472] = in_data[218975:218944] - in_data[219007:218976];
  assign out_data[109535:109504] = in_data[219039:219008] - in_data[219071:219040];
  assign out_data[109567:109536] = in_data[219103:219072] - in_data[219135:219104];
  assign out_data[109599:109568] = in_data[219167:219136] - in_data[219199:219168];
  assign out_data[109631:109600] = in_data[219231:219200] - in_data[219263:219232];
  assign out_data[109663:109632] = in_data[219295:219264] - in_data[219327:219296];
  assign out_data[109695:109664] = in_data[219359:219328] - in_data[219391:219360];
  assign out_data[109727:109696] = in_data[219423:219392] - in_data[219455:219424];
  assign out_data[10975:10944] = in_data[21919:21888] - in_data[21951:21920];
  assign out_data[109759:109728] = in_data[219487:219456] - in_data[219519:219488];
  assign out_data[109791:109760] = in_data[219551:219520] - in_data[219583:219552];
  assign out_data[109823:109792] = in_data[219615:219584] - in_data[219647:219616];
  assign out_data[109855:109824] = in_data[219679:219648] - in_data[219711:219680];
  assign out_data[109887:109856] = in_data[219743:219712] - in_data[219775:219744];
  assign out_data[109919:109888] = in_data[219807:219776] - in_data[219839:219808];
  assign out_data[109951:109920] = in_data[219871:219840] - in_data[219903:219872];
  assign out_data[109983:109952] = in_data[219935:219904] - in_data[219967:219936];
  assign out_data[110015:109984] = in_data[219999:219968] - in_data[220031:220000];
  assign out_data[110047:110016] = in_data[220063:220032] - in_data[220095:220064];
  assign out_data[11007:10976] = in_data[21983:21952] - in_data[22015:21984];
  assign out_data[110079:110048] = in_data[220127:220096] - in_data[220159:220128];
  assign out_data[110111:110080] = in_data[220191:220160] - in_data[220223:220192];
  assign out_data[110143:110112] = in_data[220255:220224] - in_data[220287:220256];
  assign out_data[110175:110144] = in_data[220319:220288] - in_data[220351:220320];
  assign out_data[110207:110176] = in_data[220383:220352] - in_data[220415:220384];
  assign out_data[110239:110208] = in_data[220447:220416] - in_data[220479:220448];
  assign out_data[110271:110240] = in_data[220511:220480] - in_data[220543:220512];
  assign out_data[110303:110272] = in_data[220575:220544] - in_data[220607:220576];
  assign out_data[110335:110304] = in_data[220639:220608] - in_data[220671:220640];
  assign out_data[110367:110336] = in_data[220703:220672] - in_data[220735:220704];
  assign out_data[11039:11008] = in_data[22047:22016] - in_data[22079:22048];
  assign out_data[110399:110368] = in_data[220767:220736] - in_data[220799:220768];
  assign out_data[110431:110400] = in_data[220831:220800] - in_data[220863:220832];
  assign out_data[110463:110432] = in_data[220895:220864] - in_data[220927:220896];
  assign out_data[110495:110464] = in_data[220959:220928] - in_data[220991:220960];
  assign out_data[110527:110496] = in_data[221023:220992] - in_data[221055:221024];
  assign out_data[110559:110528] = in_data[221087:221056] - in_data[221119:221088];
  assign out_data[110591:110560] = in_data[221151:221120] - in_data[221183:221152];
  assign out_data[110623:110592] = in_data[221215:221184] - in_data[221247:221216];
  assign out_data[110655:110624] = in_data[221279:221248] - in_data[221311:221280];
  assign out_data[110687:110656] = in_data[221343:221312] - in_data[221375:221344];
  assign out_data[11071:11040] = in_data[22111:22080] - in_data[22143:22112];
  assign out_data[110719:110688] = in_data[221407:221376] - in_data[221439:221408];
  assign out_data[110751:110720] = in_data[221471:221440] - in_data[221503:221472];
  assign out_data[110783:110752] = in_data[221535:221504] - in_data[221567:221536];
  assign out_data[110815:110784] = in_data[221599:221568] - in_data[221631:221600];
  assign out_data[110847:110816] = in_data[221663:221632] - in_data[221695:221664];
  assign out_data[110879:110848] = in_data[221727:221696] - in_data[221759:221728];
  assign out_data[110911:110880] = in_data[221791:221760] - in_data[221823:221792];
  assign out_data[110943:110912] = in_data[221855:221824] - in_data[221887:221856];
  assign out_data[110975:110944] = in_data[221919:221888] - in_data[221951:221920];
  assign out_data[111007:110976] = in_data[221983:221952] - in_data[222015:221984];
  assign out_data[11103:11072] = in_data[22175:22144] - in_data[22207:22176];
  assign out_data[111039:111008] = in_data[222047:222016] - in_data[222079:222048];
  assign out_data[111071:111040] = in_data[222111:222080] - in_data[222143:222112];
  assign out_data[111103:111072] = in_data[222175:222144] - in_data[222207:222176];
  assign out_data[111135:111104] = in_data[222239:222208] - in_data[222271:222240];
  assign out_data[111167:111136] = in_data[222303:222272] - in_data[222335:222304];
  assign out_data[111199:111168] = in_data[222367:222336] - in_data[222399:222368];
  assign out_data[111231:111200] = in_data[222431:222400] - in_data[222463:222432];
  assign out_data[111263:111232] = in_data[222495:222464] - in_data[222527:222496];
  assign out_data[111295:111264] = in_data[222559:222528] - in_data[222591:222560];
  assign out_data[111327:111296] = in_data[222623:222592] - in_data[222655:222624];
  assign out_data[11135:11104] = in_data[22239:22208] - in_data[22271:22240];
  assign out_data[111359:111328] = in_data[222687:222656] - in_data[222719:222688];
  assign out_data[111391:111360] = in_data[222751:222720] - in_data[222783:222752];
  assign out_data[111423:111392] = in_data[222815:222784] - in_data[222847:222816];
  assign out_data[111455:111424] = in_data[222879:222848] - in_data[222911:222880];
  assign out_data[111487:111456] = in_data[222943:222912] - in_data[222975:222944];
  assign out_data[111519:111488] = in_data[223007:222976] - in_data[223039:223008];
  assign out_data[111551:111520] = in_data[223071:223040] - in_data[223103:223072];
  assign out_data[111583:111552] = in_data[223135:223104] - in_data[223167:223136];
  assign out_data[111615:111584] = in_data[223199:223168] - in_data[223231:223200];
  assign out_data[111647:111616] = in_data[223263:223232] - in_data[223295:223264];
  assign out_data[11167:11136] = in_data[22303:22272] - in_data[22335:22304];
  assign out_data[111679:111648] = in_data[223327:223296] - in_data[223359:223328];
  assign out_data[111711:111680] = in_data[223391:223360] - in_data[223423:223392];
  assign out_data[111743:111712] = in_data[223455:223424] - in_data[223487:223456];
  assign out_data[111775:111744] = in_data[223519:223488] - in_data[223551:223520];
  assign out_data[111807:111776] = in_data[223583:223552] - in_data[223615:223584];
  assign out_data[111839:111808] = in_data[223647:223616] - in_data[223679:223648];
  assign out_data[111871:111840] = in_data[223711:223680] - in_data[223743:223712];
  assign out_data[111903:111872] = in_data[223775:223744] - in_data[223807:223776];
  assign out_data[111935:111904] = in_data[223839:223808] - in_data[223871:223840];
  assign out_data[111967:111936] = in_data[223903:223872] - in_data[223935:223904];
  assign out_data[1119:1088] = in_data[2207:2176] - in_data[2239:2208];
  assign out_data[11199:11168] = in_data[22367:22336] - in_data[22399:22368];
  assign out_data[111999:111968] = in_data[223967:223936] - in_data[223999:223968];
  assign out_data[112031:112000] = in_data[224031:224000] - in_data[224063:224032];
  assign out_data[112063:112032] = in_data[224095:224064] - in_data[224127:224096];
  assign out_data[112095:112064] = in_data[224159:224128] - in_data[224191:224160];
  assign out_data[112127:112096] = in_data[224223:224192] - in_data[224255:224224];
  assign out_data[112159:112128] = in_data[224287:224256] - in_data[224319:224288];
  assign out_data[112191:112160] = in_data[224351:224320] - in_data[224383:224352];
  assign out_data[112223:112192] = in_data[224415:224384] - in_data[224447:224416];
  assign out_data[112255:112224] = in_data[224479:224448] - in_data[224511:224480];
  assign out_data[112287:112256] = in_data[224543:224512] - in_data[224575:224544];
  assign out_data[11231:11200] = in_data[22431:22400] - in_data[22463:22432];
  assign out_data[112319:112288] = in_data[224607:224576] - in_data[224639:224608];
  assign out_data[112351:112320] = in_data[224671:224640] - in_data[224703:224672];
  assign out_data[112383:112352] = in_data[224735:224704] - in_data[224767:224736];
  assign out_data[112415:112384] = in_data[224799:224768] - in_data[224831:224800];
  assign out_data[112447:112416] = in_data[224863:224832] - in_data[224895:224864];
  assign out_data[112479:112448] = in_data[224927:224896] - in_data[224959:224928];
  assign out_data[112511:112480] = in_data[224991:224960] - in_data[225023:224992];
  assign out_data[112543:112512] = in_data[225055:225024] - in_data[225087:225056];
  assign out_data[112575:112544] = in_data[225119:225088] - in_data[225151:225120];
  assign out_data[112607:112576] = in_data[225183:225152] - in_data[225215:225184];
  assign out_data[11263:11232] = in_data[22495:22464] - in_data[22527:22496];
  assign out_data[112639:112608] = in_data[225247:225216] - in_data[225279:225248];
  assign out_data[112671:112640] = in_data[225311:225280] - in_data[225343:225312];
  assign out_data[112703:112672] = in_data[225375:225344] - in_data[225407:225376];
  assign out_data[112735:112704] = in_data[225439:225408] - in_data[225471:225440];
  assign out_data[112767:112736] = in_data[225503:225472] - in_data[225535:225504];
  assign out_data[112799:112768] = in_data[225567:225536] - in_data[225599:225568];
  assign out_data[112831:112800] = in_data[225631:225600] - in_data[225663:225632];
  assign out_data[112863:112832] = in_data[225695:225664] - in_data[225727:225696];
  assign out_data[112895:112864] = in_data[225759:225728] - in_data[225791:225760];
  assign out_data[112927:112896] = in_data[225823:225792] - in_data[225855:225824];
  assign out_data[11295:11264] = in_data[22559:22528] - in_data[22591:22560];
  assign out_data[112959:112928] = in_data[225887:225856] - in_data[225919:225888];
  assign out_data[112991:112960] = in_data[225951:225920] - in_data[225983:225952];
  assign out_data[113023:112992] = in_data[226015:225984] - in_data[226047:226016];
  assign out_data[113055:113024] = in_data[226079:226048] - in_data[226111:226080];
  assign out_data[113087:113056] = in_data[226143:226112] - in_data[226175:226144];
  assign out_data[113119:113088] = in_data[226207:226176] - in_data[226239:226208];
  assign out_data[113151:113120] = in_data[226271:226240] - in_data[226303:226272];
  assign out_data[113183:113152] = in_data[226335:226304] - in_data[226367:226336];
  assign out_data[113215:113184] = in_data[226399:226368] - in_data[226431:226400];
  assign out_data[113247:113216] = in_data[226463:226432] - in_data[226495:226464];
  assign out_data[11327:11296] = in_data[22623:22592] - in_data[22655:22624];
  assign out_data[113279:113248] = in_data[226527:226496] - in_data[226559:226528];
  assign out_data[113311:113280] = in_data[226591:226560] - in_data[226623:226592];
  assign out_data[113343:113312] = in_data[226655:226624] - in_data[226687:226656];
  assign out_data[113375:113344] = in_data[226719:226688] - in_data[226751:226720];
  assign out_data[113407:113376] = in_data[226783:226752] - in_data[226815:226784];
  assign out_data[113439:113408] = in_data[226847:226816] - in_data[226879:226848];
  assign out_data[113471:113440] = in_data[226911:226880] - in_data[226943:226912];
  assign out_data[113503:113472] = in_data[226975:226944] - in_data[227007:226976];
  assign out_data[113535:113504] = in_data[227039:227008] - in_data[227071:227040];
  assign out_data[113567:113536] = in_data[227103:227072] - in_data[227135:227104];
  assign out_data[11359:11328] = in_data[22687:22656] - in_data[22719:22688];
  assign out_data[113599:113568] = in_data[227167:227136] - in_data[227199:227168];
  assign out_data[113631:113600] = in_data[227231:227200] - in_data[227263:227232];
  assign out_data[113663:113632] = in_data[227295:227264] - in_data[227327:227296];
  assign out_data[113695:113664] = in_data[227359:227328] - in_data[227391:227360];
  assign out_data[113727:113696] = in_data[227423:227392] - in_data[227455:227424];
  assign out_data[113759:113728] = in_data[227487:227456] - in_data[227519:227488];
  assign out_data[113791:113760] = in_data[227551:227520] - in_data[227583:227552];
  assign out_data[113823:113792] = in_data[227615:227584] - in_data[227647:227616];
  assign out_data[113855:113824] = in_data[227679:227648] - in_data[227711:227680];
  assign out_data[113887:113856] = in_data[227743:227712] - in_data[227775:227744];
  assign out_data[11391:11360] = in_data[22751:22720] - in_data[22783:22752];
  assign out_data[113919:113888] = in_data[227807:227776] - in_data[227839:227808];
  assign out_data[113951:113920] = in_data[227871:227840] - in_data[227903:227872];
  assign out_data[113983:113952] = in_data[227935:227904] - in_data[227967:227936];
  assign out_data[114015:113984] = in_data[227999:227968] - in_data[228031:228000];
  assign out_data[114047:114016] = in_data[228063:228032] - in_data[228095:228064];
  assign out_data[114079:114048] = in_data[228127:228096] - in_data[228159:228128];
  assign out_data[114111:114080] = in_data[228191:228160] - in_data[228223:228192];
  assign out_data[114143:114112] = in_data[228255:228224] - in_data[228287:228256];
  assign out_data[114175:114144] = in_data[228319:228288] - in_data[228351:228320];
  assign out_data[114207:114176] = in_data[228383:228352] - in_data[228415:228384];
  assign out_data[11423:11392] = in_data[22815:22784] - in_data[22847:22816];
  assign out_data[114239:114208] = in_data[228447:228416] - in_data[228479:228448];
  assign out_data[114271:114240] = in_data[228511:228480] - in_data[228543:228512];
  assign out_data[114303:114272] = in_data[228575:228544] - in_data[228607:228576];
  assign out_data[114335:114304] = in_data[228639:228608] - in_data[228671:228640];
  assign out_data[114367:114336] = in_data[228703:228672] - in_data[228735:228704];
  assign out_data[114399:114368] = in_data[228767:228736] - in_data[228799:228768];
  assign out_data[114431:114400] = in_data[228831:228800] - in_data[228863:228832];
  assign out_data[114463:114432] = in_data[228895:228864] - in_data[228927:228896];
  assign out_data[114495:114464] = in_data[228959:228928] - in_data[228991:228960];
  assign out_data[114527:114496] = in_data[229023:228992] - in_data[229055:229024];
  assign out_data[11455:11424] = in_data[22879:22848] - in_data[22911:22880];
  assign out_data[114559:114528] = in_data[229087:229056] - in_data[229119:229088];
  assign out_data[114591:114560] = in_data[229151:229120] - in_data[229183:229152];
  assign out_data[114623:114592] = in_data[229215:229184] - in_data[229247:229216];
  assign out_data[114655:114624] = in_data[229279:229248] - in_data[229311:229280];
  assign out_data[114687:114656] = in_data[229343:229312] - in_data[229375:229344];
  assign out_data[114719:114688] = in_data[229407:229376] - in_data[229439:229408];
  assign out_data[114751:114720] = in_data[229471:229440] - in_data[229503:229472];
  assign out_data[114783:114752] = in_data[229535:229504] - in_data[229567:229536];
  assign out_data[114815:114784] = in_data[229599:229568] - in_data[229631:229600];
  assign out_data[114847:114816] = in_data[229663:229632] - in_data[229695:229664];
  assign out_data[11487:11456] = in_data[22943:22912] - in_data[22975:22944];
  assign out_data[114879:114848] = in_data[229727:229696] - in_data[229759:229728];
  assign out_data[114911:114880] = in_data[229791:229760] - in_data[229823:229792];
  assign out_data[114943:114912] = in_data[229855:229824] - in_data[229887:229856];
  assign out_data[114975:114944] = in_data[229919:229888] - in_data[229951:229920];
  assign out_data[115007:114976] = in_data[229983:229952] - in_data[230015:229984];
  assign out_data[115039:115008] = in_data[230047:230016] - in_data[230079:230048];
  assign out_data[115071:115040] = in_data[230111:230080] - in_data[230143:230112];
  assign out_data[115103:115072] = in_data[230175:230144] - in_data[230207:230176];
  assign out_data[115135:115104] = in_data[230239:230208] - in_data[230271:230240];
  assign out_data[115167:115136] = in_data[230303:230272] - in_data[230335:230304];
  assign out_data[1151:1120] = in_data[2271:2240] - in_data[2303:2272];
  assign out_data[11519:11488] = in_data[23007:22976] - in_data[23039:23008];
  assign out_data[115199:115168] = in_data[230367:230336] - in_data[230399:230368];
  assign out_data[115231:115200] = in_data[230431:230400] - in_data[230463:230432];
  assign out_data[115263:115232] = in_data[230495:230464] - in_data[230527:230496];
  assign out_data[115295:115264] = in_data[230559:230528] - in_data[230591:230560];
  assign out_data[115327:115296] = in_data[230623:230592] - in_data[230655:230624];
  assign out_data[115359:115328] = in_data[230687:230656] - in_data[230719:230688];
  assign out_data[115391:115360] = in_data[230751:230720] - in_data[230783:230752];
  assign out_data[115423:115392] = in_data[230815:230784] - in_data[230847:230816];
  assign out_data[115455:115424] = in_data[230879:230848] - in_data[230911:230880];
  assign out_data[115487:115456] = in_data[230943:230912] - in_data[230975:230944];
  assign out_data[11551:11520] = in_data[23071:23040] - in_data[23103:23072];
  assign out_data[115519:115488] = in_data[231007:230976] - in_data[231039:231008];
  assign out_data[115551:115520] = in_data[231071:231040] - in_data[231103:231072];
  assign out_data[115583:115552] = in_data[231135:231104] - in_data[231167:231136];
  assign out_data[115615:115584] = in_data[231199:231168] - in_data[231231:231200];
  assign out_data[115647:115616] = in_data[231263:231232] - in_data[231295:231264];
  assign out_data[115679:115648] = in_data[231327:231296] - in_data[231359:231328];
  assign out_data[115711:115680] = in_data[231391:231360] - in_data[231423:231392];
  assign out_data[115743:115712] = in_data[231455:231424] - in_data[231487:231456];
  assign out_data[115775:115744] = in_data[231519:231488] - in_data[231551:231520];
  assign out_data[115807:115776] = in_data[231583:231552] - in_data[231615:231584];
  assign out_data[11583:11552] = in_data[23135:23104] - in_data[23167:23136];
  assign out_data[115839:115808] = in_data[231647:231616] - in_data[231679:231648];
  assign out_data[115871:115840] = in_data[231711:231680] - in_data[231743:231712];
  assign out_data[115903:115872] = in_data[231775:231744] - in_data[231807:231776];
  assign out_data[115935:115904] = in_data[231839:231808] - in_data[231871:231840];
  assign out_data[115967:115936] = in_data[231903:231872] - in_data[231935:231904];
  assign out_data[115999:115968] = in_data[231967:231936] - in_data[231999:231968];
  assign out_data[116031:116000] = in_data[232031:232000] - in_data[232063:232032];
  assign out_data[116063:116032] = in_data[232095:232064] - in_data[232127:232096];
  assign out_data[116095:116064] = in_data[232159:232128] - in_data[232191:232160];
  assign out_data[116127:116096] = in_data[232223:232192] - in_data[232255:232224];
  assign out_data[11615:11584] = in_data[23199:23168] - in_data[23231:23200];
  assign out_data[116159:116128] = in_data[232287:232256] - in_data[232319:232288];
  assign out_data[116191:116160] = in_data[232351:232320] - in_data[232383:232352];
  assign out_data[116223:116192] = in_data[232415:232384] - in_data[232447:232416];
  assign out_data[116255:116224] = in_data[232479:232448] - in_data[232511:232480];
  assign out_data[116287:116256] = in_data[232543:232512] - in_data[232575:232544];
  assign out_data[116319:116288] = in_data[232607:232576] - in_data[232639:232608];
  assign out_data[116351:116320] = in_data[232671:232640] - in_data[232703:232672];
  assign out_data[116383:116352] = in_data[232735:232704] - in_data[232767:232736];
  assign out_data[116415:116384] = in_data[232799:232768] - in_data[232831:232800];
  assign out_data[116447:116416] = in_data[232863:232832] - in_data[232895:232864];
  assign out_data[11647:11616] = in_data[23263:23232] - in_data[23295:23264];
  assign out_data[116479:116448] = in_data[232927:232896] - in_data[232959:232928];
  assign out_data[116511:116480] = in_data[232991:232960] - in_data[233023:232992];
  assign out_data[116543:116512] = in_data[233055:233024] - in_data[233087:233056];
  assign out_data[116575:116544] = in_data[233119:233088] - in_data[233151:233120];
  assign out_data[116607:116576] = in_data[233183:233152] - in_data[233215:233184];
  assign out_data[116639:116608] = in_data[233247:233216] - in_data[233279:233248];
  assign out_data[116671:116640] = in_data[233311:233280] - in_data[233343:233312];
  assign out_data[116703:116672] = in_data[233375:233344] - in_data[233407:233376];
  assign out_data[116735:116704] = in_data[233439:233408] - in_data[233471:233440];
  assign out_data[116767:116736] = in_data[233503:233472] - in_data[233535:233504];
  assign out_data[11679:11648] = in_data[23327:23296] - in_data[23359:23328];
  assign out_data[116799:116768] = in_data[233567:233536] - in_data[233599:233568];
  assign out_data[116831:116800] = in_data[233631:233600] - in_data[233663:233632];
  assign out_data[116863:116832] = in_data[233695:233664] - in_data[233727:233696];
  assign out_data[116895:116864] = in_data[233759:233728] - in_data[233791:233760];
  assign out_data[116927:116896] = in_data[233823:233792] - in_data[233855:233824];
  assign out_data[116959:116928] = in_data[233887:233856] - in_data[233919:233888];
  assign out_data[116991:116960] = in_data[233951:233920] - in_data[233983:233952];
  assign out_data[117023:116992] = in_data[234015:233984] - in_data[234047:234016];
  assign out_data[117055:117024] = in_data[234079:234048] - in_data[234111:234080];
  assign out_data[117087:117056] = in_data[234143:234112] - in_data[234175:234144];
  assign out_data[11711:11680] = in_data[23391:23360] - in_data[23423:23392];
  assign out_data[117119:117088] = in_data[234207:234176] - in_data[234239:234208];
  assign out_data[117151:117120] = in_data[234271:234240] - in_data[234303:234272];
  assign out_data[117183:117152] = in_data[234335:234304] - in_data[234367:234336];
  assign out_data[117215:117184] = in_data[234399:234368] - in_data[234431:234400];
  assign out_data[117247:117216] = in_data[234463:234432] - in_data[234495:234464];
  assign out_data[117279:117248] = in_data[234527:234496] - in_data[234559:234528];
  assign out_data[117311:117280] = in_data[234591:234560] - in_data[234623:234592];
  assign out_data[117343:117312] = in_data[234655:234624] - in_data[234687:234656];
  assign out_data[117375:117344] = in_data[234719:234688] - in_data[234751:234720];
  assign out_data[117407:117376] = in_data[234783:234752] - in_data[234815:234784];
  assign out_data[11743:11712] = in_data[23455:23424] - in_data[23487:23456];
  assign out_data[117439:117408] = in_data[234847:234816] - in_data[234879:234848];
  assign out_data[117471:117440] = in_data[234911:234880] - in_data[234943:234912];
  assign out_data[117503:117472] = in_data[234975:234944] - in_data[235007:234976];
  assign out_data[117535:117504] = in_data[235039:235008] - in_data[235071:235040];
  assign out_data[117567:117536] = in_data[235103:235072] - in_data[235135:235104];
  assign out_data[117599:117568] = in_data[235167:235136] - in_data[235199:235168];
  assign out_data[117631:117600] = in_data[235231:235200] - in_data[235263:235232];
  assign out_data[117663:117632] = in_data[235295:235264] - in_data[235327:235296];
  assign out_data[117695:117664] = in_data[235359:235328] - in_data[235391:235360];
  assign out_data[117727:117696] = in_data[235423:235392] - in_data[235455:235424];
  assign out_data[11775:11744] = in_data[23519:23488] - in_data[23551:23520];
  assign out_data[117759:117728] = in_data[235487:235456] - in_data[235519:235488];
  assign out_data[117791:117760] = in_data[235551:235520] - in_data[235583:235552];
  assign out_data[117823:117792] = in_data[235615:235584] - in_data[235647:235616];
  assign out_data[117855:117824] = in_data[235679:235648] - in_data[235711:235680];
  assign out_data[117887:117856] = in_data[235743:235712] - in_data[235775:235744];
  assign out_data[117919:117888] = in_data[235807:235776] - in_data[235839:235808];
  assign out_data[117951:117920] = in_data[235871:235840] - in_data[235903:235872];
  assign out_data[117983:117952] = in_data[235935:235904] - in_data[235967:235936];
  assign out_data[118015:117984] = in_data[235999:235968] - in_data[236031:236000];
  assign out_data[118047:118016] = in_data[236063:236032] - in_data[236095:236064];
  assign out_data[11807:11776] = in_data[23583:23552] - in_data[23615:23584];
  assign out_data[118079:118048] = in_data[236127:236096] - in_data[236159:236128];
  assign out_data[118111:118080] = in_data[236191:236160] - in_data[236223:236192];
  assign out_data[118143:118112] = in_data[236255:236224] - in_data[236287:236256];
  assign out_data[118175:118144] = in_data[236319:236288] - in_data[236351:236320];
  assign out_data[118207:118176] = in_data[236383:236352] - in_data[236415:236384];
  assign out_data[118239:118208] = in_data[236447:236416] - in_data[236479:236448];
  assign out_data[118271:118240] = in_data[236511:236480] - in_data[236543:236512];
  assign out_data[118303:118272] = in_data[236575:236544] - in_data[236607:236576];
  assign out_data[118335:118304] = in_data[236639:236608] - in_data[236671:236640];
  assign out_data[118367:118336] = in_data[236703:236672] - in_data[236735:236704];
  assign out_data[1183:1152] = in_data[2335:2304] - in_data[2367:2336];
  assign out_data[11839:11808] = in_data[23647:23616] - in_data[23679:23648];
  assign out_data[118399:118368] = in_data[236767:236736] - in_data[236799:236768];
  assign out_data[118431:118400] = in_data[236831:236800] - in_data[236863:236832];
  assign out_data[118463:118432] = in_data[236895:236864] - in_data[236927:236896];
  assign out_data[118495:118464] = in_data[236959:236928] - in_data[236991:236960];
  assign out_data[118527:118496] = in_data[237023:236992] - in_data[237055:237024];
  assign out_data[118559:118528] = in_data[237087:237056] - in_data[237119:237088];
  assign out_data[118591:118560] = in_data[237151:237120] - in_data[237183:237152];
  assign out_data[118623:118592] = in_data[237215:237184] - in_data[237247:237216];
  assign out_data[118655:118624] = in_data[237279:237248] - in_data[237311:237280];
  assign out_data[118687:118656] = in_data[237343:237312] - in_data[237375:237344];
  assign out_data[11871:11840] = in_data[23711:23680] - in_data[23743:23712];
  assign out_data[118719:118688] = in_data[237407:237376] - in_data[237439:237408];
  assign out_data[118751:118720] = in_data[237471:237440] - in_data[237503:237472];
  assign out_data[118783:118752] = in_data[237535:237504] - in_data[237567:237536];
  assign out_data[118815:118784] = in_data[237599:237568] - in_data[237631:237600];
  assign out_data[118847:118816] = in_data[237663:237632] - in_data[237695:237664];
  assign out_data[118879:118848] = in_data[237727:237696] - in_data[237759:237728];
  assign out_data[118911:118880] = in_data[237791:237760] - in_data[237823:237792];
  assign out_data[118943:118912] = in_data[237855:237824] - in_data[237887:237856];
  assign out_data[118975:118944] = in_data[237919:237888] - in_data[237951:237920];
  assign out_data[119007:118976] = in_data[237983:237952] - in_data[238015:237984];
  assign out_data[11903:11872] = in_data[23775:23744] - in_data[23807:23776];
  assign out_data[119039:119008] = in_data[238047:238016] - in_data[238079:238048];
  assign out_data[119071:119040] = in_data[238111:238080] - in_data[238143:238112];
  assign out_data[119103:119072] = in_data[238175:238144] - in_data[238207:238176];
  assign out_data[119135:119104] = in_data[238239:238208] - in_data[238271:238240];
  assign out_data[119167:119136] = in_data[238303:238272] - in_data[238335:238304];
  assign out_data[119199:119168] = in_data[238367:238336] - in_data[238399:238368];
  assign out_data[119231:119200] = in_data[238431:238400] - in_data[238463:238432];
  assign out_data[119263:119232] = in_data[238495:238464] - in_data[238527:238496];
  assign out_data[119295:119264] = in_data[238559:238528] - in_data[238591:238560];
  assign out_data[119327:119296] = in_data[238623:238592] - in_data[238655:238624];
  assign out_data[11935:11904] = in_data[23839:23808] - in_data[23871:23840];
  assign out_data[119359:119328] = in_data[238687:238656] - in_data[238719:238688];
  assign out_data[119391:119360] = in_data[238751:238720] - in_data[238783:238752];
  assign out_data[119423:119392] = in_data[238815:238784] - in_data[238847:238816];
  assign out_data[119455:119424] = in_data[238879:238848] - in_data[238911:238880];
  assign out_data[119487:119456] = in_data[238943:238912] - in_data[238975:238944];
  assign out_data[119519:119488] = in_data[239007:238976] - in_data[239039:239008];
  assign out_data[119551:119520] = in_data[239071:239040] - in_data[239103:239072];
  assign out_data[119583:119552] = in_data[239135:239104] - in_data[239167:239136];
  assign out_data[119615:119584] = in_data[239199:239168] - in_data[239231:239200];
  assign out_data[119647:119616] = in_data[239263:239232] - in_data[239295:239264];
  assign out_data[11967:11936] = in_data[23903:23872] - in_data[23935:23904];
  assign out_data[119679:119648] = in_data[239327:239296] - in_data[239359:239328];
  assign out_data[119711:119680] = in_data[239391:239360] - in_data[239423:239392];
  assign out_data[119743:119712] = in_data[239455:239424] - in_data[239487:239456];
  assign out_data[119775:119744] = in_data[239519:239488] - in_data[239551:239520];
  assign out_data[119807:119776] = in_data[239583:239552] - in_data[239615:239584];
  assign out_data[119839:119808] = in_data[239647:239616] - in_data[239679:239648];
  assign out_data[119871:119840] = in_data[239711:239680] - in_data[239743:239712];
  assign out_data[119903:119872] = in_data[239775:239744] - in_data[239807:239776];
  assign out_data[119935:119904] = in_data[239839:239808] - in_data[239871:239840];
  assign out_data[119967:119936] = in_data[239903:239872] - in_data[239935:239904];
  assign out_data[11999:11968] = in_data[23967:23936] - in_data[23999:23968];
  assign out_data[119999:119968] = in_data[239967:239936] - in_data[239999:239968];
  assign out_data[120031:120000] = in_data[240031:240000] - in_data[240063:240032];
  assign out_data[120063:120032] = in_data[240095:240064] - in_data[240127:240096];
  assign out_data[120095:120064] = in_data[240159:240128] - in_data[240191:240160];
  assign out_data[120127:120096] = in_data[240223:240192] - in_data[240255:240224];
  assign out_data[120159:120128] = in_data[240287:240256] - in_data[240319:240288];
  assign out_data[120191:120160] = in_data[240351:240320] - in_data[240383:240352];
  assign out_data[120223:120192] = in_data[240415:240384] - in_data[240447:240416];
  assign out_data[120255:120224] = in_data[240479:240448] - in_data[240511:240480];
  assign out_data[120287:120256] = in_data[240543:240512] - in_data[240575:240544];
  assign out_data[12031:12000] = in_data[24031:24000] - in_data[24063:24032];
  assign out_data[120319:120288] = in_data[240607:240576] - in_data[240639:240608];
  assign out_data[120351:120320] = in_data[240671:240640] - in_data[240703:240672];
  assign out_data[120383:120352] = in_data[240735:240704] - in_data[240767:240736];
  assign out_data[120415:120384] = in_data[240799:240768] - in_data[240831:240800];
  assign out_data[120447:120416] = in_data[240863:240832] - in_data[240895:240864];
  assign out_data[120479:120448] = in_data[240927:240896] - in_data[240959:240928];
  assign out_data[120511:120480] = in_data[240991:240960] - in_data[241023:240992];
  assign out_data[120543:120512] = in_data[241055:241024] - in_data[241087:241056];
  assign out_data[120575:120544] = in_data[241119:241088] - in_data[241151:241120];
  assign out_data[120607:120576] = in_data[241183:241152] - in_data[241215:241184];
  assign out_data[12063:12032] = in_data[24095:24064] - in_data[24127:24096];
  assign out_data[120639:120608] = in_data[241247:241216] - in_data[241279:241248];
  assign out_data[120671:120640] = in_data[241311:241280] - in_data[241343:241312];
  assign out_data[120703:120672] = in_data[241375:241344] - in_data[241407:241376];
  assign out_data[120735:120704] = in_data[241439:241408] - in_data[241471:241440];
  assign out_data[120767:120736] = in_data[241503:241472] - in_data[241535:241504];
  assign out_data[120799:120768] = in_data[241567:241536] - in_data[241599:241568];
  assign out_data[120831:120800] = in_data[241631:241600] - in_data[241663:241632];
  assign out_data[120863:120832] = in_data[241695:241664] - in_data[241727:241696];
  assign out_data[120895:120864] = in_data[241759:241728] - in_data[241791:241760];
  assign out_data[120927:120896] = in_data[241823:241792] - in_data[241855:241824];
  assign out_data[12095:12064] = in_data[24159:24128] - in_data[24191:24160];
  assign out_data[120959:120928] = in_data[241887:241856] - in_data[241919:241888];
  assign out_data[120991:120960] = in_data[241951:241920] - in_data[241983:241952];
  assign out_data[121023:120992] = in_data[242015:241984] - in_data[242047:242016];
  assign out_data[121055:121024] = in_data[242079:242048] - in_data[242111:242080];
  assign out_data[121087:121056] = in_data[242143:242112] - in_data[242175:242144];
  assign out_data[121119:121088] = in_data[242207:242176] - in_data[242239:242208];
  assign out_data[121151:121120] = in_data[242271:242240] - in_data[242303:242272];
  assign out_data[121183:121152] = in_data[242335:242304] - in_data[242367:242336];
  assign out_data[121215:121184] = in_data[242399:242368] - in_data[242431:242400];
  assign out_data[121247:121216] = in_data[242463:242432] - in_data[242495:242464];
  assign out_data[12127:12096] = in_data[24223:24192] - in_data[24255:24224];
  assign out_data[121279:121248] = in_data[242527:242496] - in_data[242559:242528];
  assign out_data[121311:121280] = in_data[242591:242560] - in_data[242623:242592];
  assign out_data[121343:121312] = in_data[242655:242624] - in_data[242687:242656];
  assign out_data[121375:121344] = in_data[242719:242688] - in_data[242751:242720];
  assign out_data[121407:121376] = in_data[242783:242752] - in_data[242815:242784];
  assign out_data[121439:121408] = in_data[242847:242816] - in_data[242879:242848];
  assign out_data[121471:121440] = in_data[242911:242880] - in_data[242943:242912];
  assign out_data[121503:121472] = in_data[242975:242944] - in_data[243007:242976];
  assign out_data[121535:121504] = in_data[243039:243008] - in_data[243071:243040];
  assign out_data[121567:121536] = in_data[243103:243072] - in_data[243135:243104];
  assign out_data[1215:1184] = in_data[2399:2368] - in_data[2431:2400];
  assign out_data[12159:12128] = in_data[24287:24256] - in_data[24319:24288];
  assign out_data[121599:121568] = in_data[243167:243136] - in_data[243199:243168];
  assign out_data[121631:121600] = in_data[243231:243200] - in_data[243263:243232];
  assign out_data[121663:121632] = in_data[243295:243264] - in_data[243327:243296];
  assign out_data[121695:121664] = in_data[243359:243328] - in_data[243391:243360];
  assign out_data[121727:121696] = in_data[243423:243392] - in_data[243455:243424];
  assign out_data[121759:121728] = in_data[243487:243456] - in_data[243519:243488];
  assign out_data[121791:121760] = in_data[243551:243520] - in_data[243583:243552];
  assign out_data[121823:121792] = in_data[243615:243584] - in_data[243647:243616];
  assign out_data[121855:121824] = in_data[243679:243648] - in_data[243711:243680];
  assign out_data[121887:121856] = in_data[243743:243712] - in_data[243775:243744];
  assign out_data[12191:12160] = in_data[24351:24320] - in_data[24383:24352];
  assign out_data[121919:121888] = in_data[243807:243776] - in_data[243839:243808];
  assign out_data[121951:121920] = in_data[243871:243840] - in_data[243903:243872];
  assign out_data[121983:121952] = in_data[243935:243904] - in_data[243967:243936];
  assign out_data[122015:121984] = in_data[243999:243968] - in_data[244031:244000];
  assign out_data[122047:122016] = in_data[244063:244032] - in_data[244095:244064];
  assign out_data[122079:122048] = in_data[244127:244096] - in_data[244159:244128];
  assign out_data[122111:122080] = in_data[244191:244160] - in_data[244223:244192];
  assign out_data[122143:122112] = in_data[244255:244224] - in_data[244287:244256];
  assign out_data[122175:122144] = in_data[244319:244288] - in_data[244351:244320];
  assign out_data[122207:122176] = in_data[244383:244352] - in_data[244415:244384];
  assign out_data[12223:12192] = in_data[24415:24384] - in_data[24447:24416];
  assign out_data[122239:122208] = in_data[244447:244416] - in_data[244479:244448];
  assign out_data[122271:122240] = in_data[244511:244480] - in_data[244543:244512];
  assign out_data[122303:122272] = in_data[244575:244544] - in_data[244607:244576];
  assign out_data[122335:122304] = in_data[244639:244608] - in_data[244671:244640];
  assign out_data[122367:122336] = in_data[244703:244672] - in_data[244735:244704];
  assign out_data[122399:122368] = in_data[244767:244736] - in_data[244799:244768];
  assign out_data[122431:122400] = in_data[244831:244800] - in_data[244863:244832];
  assign out_data[122463:122432] = in_data[244895:244864] - in_data[244927:244896];
  assign out_data[122495:122464] = in_data[244959:244928] - in_data[244991:244960];
  assign out_data[122527:122496] = in_data[245023:244992] - in_data[245055:245024];
  assign out_data[12255:12224] = in_data[24479:24448] - in_data[24511:24480];
  assign out_data[122559:122528] = in_data[245087:245056] - in_data[245119:245088];
  assign out_data[122591:122560] = in_data[245151:245120] - in_data[245183:245152];
  assign out_data[122623:122592] = in_data[245215:245184] - in_data[245247:245216];
  assign out_data[122655:122624] = in_data[245279:245248] - in_data[245311:245280];
  assign out_data[122687:122656] = in_data[245343:245312] - in_data[245375:245344];
  assign out_data[122719:122688] = in_data[245407:245376] - in_data[245439:245408];
  assign out_data[122751:122720] = in_data[245471:245440] - in_data[245503:245472];
  assign out_data[122783:122752] = in_data[245535:245504] - in_data[245567:245536];
  assign out_data[122815:122784] = in_data[245599:245568] - in_data[245631:245600];
  assign out_data[122847:122816] = in_data[245663:245632] - in_data[245695:245664];
  assign out_data[12287:12256] = in_data[24543:24512] - in_data[24575:24544];
  assign out_data[122879:122848] = in_data[245727:245696] - in_data[245759:245728];
  assign out_data[122911:122880] = in_data[245791:245760] - in_data[245823:245792];
  assign out_data[122943:122912] = in_data[245855:245824] - in_data[245887:245856];
  assign out_data[122975:122944] = in_data[245919:245888] - in_data[245951:245920];
  assign out_data[123007:122976] = in_data[245983:245952] - in_data[246015:245984];
  assign out_data[123039:123008] = in_data[246047:246016] - in_data[246079:246048];
  assign out_data[123071:123040] = in_data[246111:246080] - in_data[246143:246112];
  assign out_data[123103:123072] = in_data[246175:246144] - in_data[246207:246176];
  assign out_data[123135:123104] = in_data[246239:246208] - in_data[246271:246240];
  assign out_data[123167:123136] = in_data[246303:246272] - in_data[246335:246304];
  assign out_data[12319:12288] = in_data[24607:24576] - in_data[24639:24608];
  assign out_data[123199:123168] = in_data[246367:246336] - in_data[246399:246368];
  assign out_data[123231:123200] = in_data[246431:246400] - in_data[246463:246432];
  assign out_data[123263:123232] = in_data[246495:246464] - in_data[246527:246496];
  assign out_data[123295:123264] = in_data[246559:246528] - in_data[246591:246560];
  assign out_data[123327:123296] = in_data[246623:246592] - in_data[246655:246624];
  assign out_data[123359:123328] = in_data[246687:246656] - in_data[246719:246688];
  assign out_data[123391:123360] = in_data[246751:246720] - in_data[246783:246752];
  assign out_data[123423:123392] = in_data[246815:246784] - in_data[246847:246816];
  assign out_data[123455:123424] = in_data[246879:246848] - in_data[246911:246880];
  assign out_data[123487:123456] = in_data[246943:246912] - in_data[246975:246944];
  assign out_data[12351:12320] = in_data[24671:24640] - in_data[24703:24672];
  assign out_data[123519:123488] = in_data[247007:246976] - in_data[247039:247008];
  assign out_data[123551:123520] = in_data[247071:247040] - in_data[247103:247072];
  assign out_data[123583:123552] = in_data[247135:247104] - in_data[247167:247136];
  assign out_data[123615:123584] = in_data[247199:247168] - in_data[247231:247200];
  assign out_data[123647:123616] = in_data[247263:247232] - in_data[247295:247264];
  assign out_data[123679:123648] = in_data[247327:247296] - in_data[247359:247328];
  assign out_data[123711:123680] = in_data[247391:247360] - in_data[247423:247392];
  assign out_data[123743:123712] = in_data[247455:247424] - in_data[247487:247456];
  assign out_data[123775:123744] = in_data[247519:247488] - in_data[247551:247520];
  assign out_data[123807:123776] = in_data[247583:247552] - in_data[247615:247584];
  assign out_data[12383:12352] = in_data[24735:24704] - in_data[24767:24736];
  assign out_data[123839:123808] = in_data[247647:247616] - in_data[247679:247648];
  assign out_data[123871:123840] = in_data[247711:247680] - in_data[247743:247712];
  assign out_data[123903:123872] = in_data[247775:247744] - in_data[247807:247776];
  assign out_data[123935:123904] = in_data[247839:247808] - in_data[247871:247840];
  assign out_data[123967:123936] = in_data[247903:247872] - in_data[247935:247904];
  assign out_data[123999:123968] = in_data[247967:247936] - in_data[247999:247968];
  assign out_data[124031:124000] = in_data[248031:248000] - in_data[248063:248032];
  assign out_data[124063:124032] = in_data[248095:248064] - in_data[248127:248096];
  assign out_data[124095:124064] = in_data[248159:248128] - in_data[248191:248160];
  assign out_data[124127:124096] = in_data[248223:248192] - in_data[248255:248224];
  assign out_data[12415:12384] = in_data[24799:24768] - in_data[24831:24800];
  assign out_data[124159:124128] = in_data[248287:248256] - in_data[248319:248288];
  assign out_data[124191:124160] = in_data[248351:248320] - in_data[248383:248352];
  assign out_data[124223:124192] = in_data[248415:248384] - in_data[248447:248416];
  assign out_data[124255:124224] = in_data[248479:248448] - in_data[248511:248480];
  assign out_data[124287:124256] = in_data[248543:248512] - in_data[248575:248544];
  assign out_data[124319:124288] = in_data[248607:248576] - in_data[248639:248608];
  assign out_data[124351:124320] = in_data[248671:248640] - in_data[248703:248672];
  assign out_data[124383:124352] = in_data[248735:248704] - in_data[248767:248736];
  assign out_data[124415:124384] = in_data[248799:248768] - in_data[248831:248800];
  assign out_data[124447:124416] = in_data[248863:248832] - in_data[248895:248864];
  assign out_data[12447:12416] = in_data[24863:24832] - in_data[24895:24864];
  assign out_data[124479:124448] = in_data[248927:248896] - in_data[248959:248928];
  assign out_data[124511:124480] = in_data[248991:248960] - in_data[249023:248992];
  assign out_data[124543:124512] = in_data[249055:249024] - in_data[249087:249056];
  assign out_data[124575:124544] = in_data[249119:249088] - in_data[249151:249120];
  assign out_data[124607:124576] = in_data[249183:249152] - in_data[249215:249184];
  assign out_data[124639:124608] = in_data[249247:249216] - in_data[249279:249248];
  assign out_data[124671:124640] = in_data[249311:249280] - in_data[249343:249312];
  assign out_data[124703:124672] = in_data[249375:249344] - in_data[249407:249376];
  assign out_data[124735:124704] = in_data[249439:249408] - in_data[249471:249440];
  assign out_data[124767:124736] = in_data[249503:249472] - in_data[249535:249504];
  assign out_data[1247:1216] = in_data[2463:2432] - in_data[2495:2464];
  assign out_data[12479:12448] = in_data[24927:24896] - in_data[24959:24928];
  assign out_data[124799:124768] = in_data[249567:249536] - in_data[249599:249568];
  assign out_data[124831:124800] = in_data[249631:249600] - in_data[249663:249632];
  assign out_data[124863:124832] = in_data[249695:249664] - in_data[249727:249696];
  assign out_data[124895:124864] = in_data[249759:249728] - in_data[249791:249760];
  assign out_data[124927:124896] = in_data[249823:249792] - in_data[249855:249824];
  assign out_data[124959:124928] = in_data[249887:249856] - in_data[249919:249888];
  assign out_data[124991:124960] = in_data[249951:249920] - in_data[249983:249952];
  assign out_data[125023:124992] = in_data[250015:249984] - in_data[250047:250016];
  assign out_data[125055:125024] = in_data[250079:250048] - in_data[250111:250080];
  assign out_data[125087:125056] = in_data[250143:250112] - in_data[250175:250144];
  assign out_data[12511:12480] = in_data[24991:24960] - in_data[25023:24992];
  assign out_data[125119:125088] = in_data[250207:250176] - in_data[250239:250208];
  assign out_data[125151:125120] = in_data[250271:250240] - in_data[250303:250272];
  assign out_data[125183:125152] = in_data[250335:250304] - in_data[250367:250336];
  assign out_data[125215:125184] = in_data[250399:250368] - in_data[250431:250400];
  assign out_data[125247:125216] = in_data[250463:250432] - in_data[250495:250464];
  assign out_data[125279:125248] = in_data[250527:250496] - in_data[250559:250528];
  assign out_data[125311:125280] = in_data[250591:250560] - in_data[250623:250592];
  assign out_data[125343:125312] = in_data[250655:250624] - in_data[250687:250656];
  assign out_data[125375:125344] = in_data[250719:250688] - in_data[250751:250720];
  assign out_data[125407:125376] = in_data[250783:250752] - in_data[250815:250784];
  assign out_data[12543:12512] = in_data[25055:25024] - in_data[25087:25056];
  assign out_data[125439:125408] = in_data[250847:250816] - in_data[250879:250848];
  assign out_data[125471:125440] = in_data[250911:250880] - in_data[250943:250912];
  assign out_data[125503:125472] = in_data[250975:250944] - in_data[251007:250976];
  assign out_data[125535:125504] = in_data[251039:251008] - in_data[251071:251040];
  assign out_data[125567:125536] = in_data[251103:251072] - in_data[251135:251104];
  assign out_data[125599:125568] = in_data[251167:251136] - in_data[251199:251168];
  assign out_data[125631:125600] = in_data[251231:251200] - in_data[251263:251232];
  assign out_data[125663:125632] = in_data[251295:251264] - in_data[251327:251296];
  assign out_data[125695:125664] = in_data[251359:251328] - in_data[251391:251360];
  assign out_data[125727:125696] = in_data[251423:251392] - in_data[251455:251424];
  assign out_data[12575:12544] = in_data[25119:25088] - in_data[25151:25120];
  assign out_data[125759:125728] = in_data[251487:251456] - in_data[251519:251488];
  assign out_data[125791:125760] = in_data[251551:251520] - in_data[251583:251552];
  assign out_data[125823:125792] = in_data[251615:251584] - in_data[251647:251616];
  assign out_data[125855:125824] = in_data[251679:251648] - in_data[251711:251680];
  assign out_data[125887:125856] = in_data[251743:251712] - in_data[251775:251744];
  assign out_data[125919:125888] = in_data[251807:251776] - in_data[251839:251808];
  assign out_data[125951:125920] = in_data[251871:251840] - in_data[251903:251872];
  assign out_data[125983:125952] = in_data[251935:251904] - in_data[251967:251936];
  assign out_data[126015:125984] = in_data[251999:251968] - in_data[252031:252000];
  assign out_data[126047:126016] = in_data[252063:252032] - in_data[252095:252064];
  assign out_data[12607:12576] = in_data[25183:25152] - in_data[25215:25184];
  assign out_data[126079:126048] = in_data[252127:252096] - in_data[252159:252128];
  assign out_data[126111:126080] = in_data[252191:252160] - in_data[252223:252192];
  assign out_data[126143:126112] = in_data[252255:252224] - in_data[252287:252256];
  assign out_data[126175:126144] = in_data[252319:252288] - in_data[252351:252320];
  assign out_data[126207:126176] = in_data[252383:252352] - in_data[252415:252384];
  assign out_data[126239:126208] = in_data[252447:252416] - in_data[252479:252448];
  assign out_data[126271:126240] = in_data[252511:252480] - in_data[252543:252512];
  assign out_data[126303:126272] = in_data[252575:252544] - in_data[252607:252576];
  assign out_data[126335:126304] = in_data[252639:252608] - in_data[252671:252640];
  assign out_data[126367:126336] = in_data[252703:252672] - in_data[252735:252704];
  assign out_data[12639:12608] = in_data[25247:25216] - in_data[25279:25248];
  assign out_data[126399:126368] = in_data[252767:252736] - in_data[252799:252768];
  assign out_data[126431:126400] = in_data[252831:252800] - in_data[252863:252832];
  assign out_data[126463:126432] = in_data[252895:252864] - in_data[252927:252896];
  assign out_data[126495:126464] = in_data[252959:252928] - in_data[252991:252960];
  assign out_data[126527:126496] = in_data[253023:252992] - in_data[253055:253024];
  assign out_data[126559:126528] = in_data[253087:253056] - in_data[253119:253088];
  assign out_data[126591:126560] = in_data[253151:253120] - in_data[253183:253152];
  assign out_data[126623:126592] = in_data[253215:253184] - in_data[253247:253216];
  assign out_data[126655:126624] = in_data[253279:253248] - in_data[253311:253280];
  assign out_data[126687:126656] = in_data[253343:253312] - in_data[253375:253344];
  assign out_data[12671:12640] = in_data[25311:25280] - in_data[25343:25312];
  assign out_data[126719:126688] = in_data[253407:253376] - in_data[253439:253408];
  assign out_data[126751:126720] = in_data[253471:253440] - in_data[253503:253472];
  assign out_data[126783:126752] = in_data[253535:253504] - in_data[253567:253536];
  assign out_data[126815:126784] = in_data[253599:253568] - in_data[253631:253600];
  assign out_data[126847:126816] = in_data[253663:253632] - in_data[253695:253664];
  assign out_data[126879:126848] = in_data[253727:253696] - in_data[253759:253728];
  assign out_data[126911:126880] = in_data[253791:253760] - in_data[253823:253792];
  assign out_data[126943:126912] = in_data[253855:253824] - in_data[253887:253856];
  assign out_data[126975:126944] = in_data[253919:253888] - in_data[253951:253920];
  assign out_data[127007:126976] = in_data[253983:253952] - in_data[254015:253984];
  assign out_data[12703:12672] = in_data[25375:25344] - in_data[25407:25376];
  assign out_data[127039:127008] = in_data[254047:254016] - in_data[254079:254048];
  assign out_data[127071:127040] = in_data[254111:254080] - in_data[254143:254112];
  assign out_data[127103:127072] = in_data[254175:254144] - in_data[254207:254176];
  assign out_data[127135:127104] = in_data[254239:254208] - in_data[254271:254240];
  assign out_data[127167:127136] = in_data[254303:254272] - in_data[254335:254304];
  assign out_data[127199:127168] = in_data[254367:254336] - in_data[254399:254368];
  assign out_data[127231:127200] = in_data[254431:254400] - in_data[254463:254432];
  assign out_data[127263:127232] = in_data[254495:254464] - in_data[254527:254496];
  assign out_data[127295:127264] = in_data[254559:254528] - in_data[254591:254560];
  assign out_data[127327:127296] = in_data[254623:254592] - in_data[254655:254624];
  assign out_data[12735:12704] = in_data[25439:25408] - in_data[25471:25440];
  assign out_data[127359:127328] = in_data[254687:254656] - in_data[254719:254688];
  assign out_data[127391:127360] = in_data[254751:254720] - in_data[254783:254752];
  assign out_data[127423:127392] = in_data[254815:254784] - in_data[254847:254816];
  assign out_data[127455:127424] = in_data[254879:254848] - in_data[254911:254880];
  assign out_data[127487:127456] = in_data[254943:254912] - in_data[254975:254944];
  assign out_data[127519:127488] = in_data[255007:254976] - in_data[255039:255008];
  assign out_data[127551:127520] = in_data[255071:255040] - in_data[255103:255072];
  assign out_data[127583:127552] = in_data[255135:255104] - in_data[255167:255136];
  assign out_data[127615:127584] = in_data[255199:255168] - in_data[255231:255200];
  assign out_data[127647:127616] = in_data[255263:255232] - in_data[255295:255264];
  assign out_data[12767:12736] = in_data[25503:25472] - in_data[25535:25504];
  assign out_data[127679:127648] = in_data[255327:255296] - in_data[255359:255328];
  assign out_data[127711:127680] = in_data[255391:255360] - in_data[255423:255392];
  assign out_data[127743:127712] = in_data[255455:255424] - in_data[255487:255456];
  assign out_data[127775:127744] = in_data[255519:255488] - in_data[255551:255520];
  assign out_data[127807:127776] = in_data[255583:255552] - in_data[255615:255584];
  assign out_data[127839:127808] = in_data[255647:255616] - in_data[255679:255648];
  assign out_data[127871:127840] = in_data[255711:255680] - in_data[255743:255712];
  assign out_data[127903:127872] = in_data[255775:255744] - in_data[255807:255776];
  assign out_data[127935:127904] = in_data[255839:255808] - in_data[255871:255840];
  assign out_data[127967:127936] = in_data[255903:255872] - in_data[255935:255904];
  assign out_data[127:96] = in_data[223:192] - in_data[255:224];
  assign out_data[1279:1248] = in_data[2527:2496] - in_data[2559:2528];
  assign out_data[12799:12768] = in_data[25567:25536] - in_data[25599:25568];
  assign out_data[127999:127968] = in_data[255967:255936] - in_data[255999:255968];
  assign out_data[128031:128000] = in_data[256031:256000] - in_data[256063:256032];
  assign out_data[128063:128032] = in_data[256095:256064] - in_data[256127:256096];
  assign out_data[128095:128064] = in_data[256159:256128] - in_data[256191:256160];
  assign out_data[128127:128096] = in_data[256223:256192] - in_data[256255:256224];
  assign out_data[128159:128128] = in_data[256287:256256] - in_data[256319:256288];
  assign out_data[128191:128160] = in_data[256351:256320] - in_data[256383:256352];
  assign out_data[128223:128192] = in_data[256415:256384] - in_data[256447:256416];
  assign out_data[128255:128224] = in_data[256479:256448] - in_data[256511:256480];
  assign out_data[128287:128256] = in_data[256543:256512] - in_data[256575:256544];
  assign out_data[12831:12800] = in_data[25631:25600] - in_data[25663:25632];
  assign out_data[128319:128288] = in_data[256607:256576] - in_data[256639:256608];
  assign out_data[128351:128320] = in_data[256671:256640] - in_data[256703:256672];
  assign out_data[128383:128352] = in_data[256735:256704] - in_data[256767:256736];
  assign out_data[128415:128384] = in_data[256799:256768] - in_data[256831:256800];
  assign out_data[128447:128416] = in_data[256863:256832] - in_data[256895:256864];
  assign out_data[128479:128448] = in_data[256927:256896] - in_data[256959:256928];
  assign out_data[128511:128480] = in_data[256991:256960] - in_data[257023:256992];
  assign out_data[128543:128512] = in_data[257055:257024] - in_data[257087:257056];
  assign out_data[128575:128544] = in_data[257119:257088] - in_data[257151:257120];
  assign out_data[128607:128576] = in_data[257183:257152] - in_data[257215:257184];
  assign out_data[12863:12832] = in_data[25695:25664] - in_data[25727:25696];
  assign out_data[128639:128608] = in_data[257247:257216] - in_data[257279:257248];
  assign out_data[128671:128640] = in_data[257311:257280] - in_data[257343:257312];
  assign out_data[128703:128672] = in_data[257375:257344] - in_data[257407:257376];
  assign out_data[128735:128704] = in_data[257439:257408] - in_data[257471:257440];
  assign out_data[128767:128736] = in_data[257503:257472] - in_data[257535:257504];
  assign out_data[128799:128768] = in_data[257567:257536] - in_data[257599:257568];
  assign out_data[128831:128800] = in_data[257631:257600] - in_data[257663:257632];
  assign out_data[128863:128832] = in_data[257695:257664] - in_data[257727:257696];
  assign out_data[128895:128864] = in_data[257759:257728] - in_data[257791:257760];
  assign out_data[128927:128896] = in_data[257823:257792] - in_data[257855:257824];
  assign out_data[12895:12864] = in_data[25759:25728] - in_data[25791:25760];
  assign out_data[128959:128928] = in_data[257887:257856] - in_data[257919:257888];
  assign out_data[128991:128960] = in_data[257951:257920] - in_data[257983:257952];
  assign out_data[129023:128992] = in_data[258015:257984] - in_data[258047:258016];
  assign out_data[129055:129024] = in_data[258079:258048] - in_data[258111:258080];
  assign out_data[129087:129056] = in_data[258143:258112] - in_data[258175:258144];
  assign out_data[129119:129088] = in_data[258207:258176] - in_data[258239:258208];
  assign out_data[129151:129120] = in_data[258271:258240] - in_data[258303:258272];
  assign out_data[129183:129152] = in_data[258335:258304] - in_data[258367:258336];
  assign out_data[129215:129184] = in_data[258399:258368] - in_data[258431:258400];
  assign out_data[129247:129216] = in_data[258463:258432] - in_data[258495:258464];
  assign out_data[12927:12896] = in_data[25823:25792] - in_data[25855:25824];
  assign out_data[129279:129248] = in_data[258527:258496] - in_data[258559:258528];
  assign out_data[129311:129280] = in_data[258591:258560] - in_data[258623:258592];
  assign out_data[129343:129312] = in_data[258655:258624] - in_data[258687:258656];
  assign out_data[129375:129344] = in_data[258719:258688] - in_data[258751:258720];
  assign out_data[129407:129376] = in_data[258783:258752] - in_data[258815:258784];
  assign out_data[129439:129408] = in_data[258847:258816] - in_data[258879:258848];
  assign out_data[129471:129440] = in_data[258911:258880] - in_data[258943:258912];
  assign out_data[129503:129472] = in_data[258975:258944] - in_data[259007:258976];
  assign out_data[129535:129504] = in_data[259039:259008] - in_data[259071:259040];
  assign out_data[129567:129536] = in_data[259103:259072] - in_data[259135:259104];
  assign out_data[12959:12928] = in_data[25887:25856] - in_data[25919:25888];
  assign out_data[129599:129568] = in_data[259167:259136] - in_data[259199:259168];
  assign out_data[129631:129600] = in_data[259231:259200] - in_data[259263:259232];
  assign out_data[129663:129632] = in_data[259295:259264] - in_data[259327:259296];
  assign out_data[129695:129664] = in_data[259359:259328] - in_data[259391:259360];
  assign out_data[129727:129696] = in_data[259423:259392] - in_data[259455:259424];
  assign out_data[129759:129728] = in_data[259487:259456] - in_data[259519:259488];
  assign out_data[129791:129760] = in_data[259551:259520] - in_data[259583:259552];
  assign out_data[129823:129792] = in_data[259615:259584] - in_data[259647:259616];
  assign out_data[129855:129824] = in_data[259679:259648] - in_data[259711:259680];
  assign out_data[129887:129856] = in_data[259743:259712] - in_data[259775:259744];
  assign out_data[12991:12960] = in_data[25951:25920] - in_data[25983:25952];
  assign out_data[129919:129888] = in_data[259807:259776] - in_data[259839:259808];
  assign out_data[129951:129920] = in_data[259871:259840] - in_data[259903:259872];
  assign out_data[129983:129952] = in_data[259935:259904] - in_data[259967:259936];
  assign out_data[130015:129984] = in_data[259999:259968] - in_data[260031:260000];
  assign out_data[130047:130016] = in_data[260063:260032] - in_data[260095:260064];
  assign out_data[130079:130048] = in_data[260127:260096] - in_data[260159:260128];
  assign out_data[130111:130080] = in_data[260191:260160] - in_data[260223:260192];
  assign out_data[130143:130112] = in_data[260255:260224] - in_data[260287:260256];
  assign out_data[130175:130144] = in_data[260319:260288] - in_data[260351:260320];
  assign out_data[130207:130176] = in_data[260383:260352] - in_data[260415:260384];
  assign out_data[13023:12992] = in_data[26015:25984] - in_data[26047:26016];
  assign out_data[130239:130208] = in_data[260447:260416] - in_data[260479:260448];
  assign out_data[130271:130240] = in_data[260511:260480] - in_data[260543:260512];
  assign out_data[130303:130272] = in_data[260575:260544] - in_data[260607:260576];
  assign out_data[130335:130304] = in_data[260639:260608] - in_data[260671:260640];
  assign out_data[130367:130336] = in_data[260703:260672] - in_data[260735:260704];
  assign out_data[130399:130368] = in_data[260767:260736] - in_data[260799:260768];
  assign out_data[130431:130400] = in_data[260831:260800] - in_data[260863:260832];
  assign out_data[130463:130432] = in_data[260895:260864] - in_data[260927:260896];
  assign out_data[130495:130464] = in_data[260959:260928] - in_data[260991:260960];
  assign out_data[130527:130496] = in_data[261023:260992] - in_data[261055:261024];
  assign out_data[13055:13024] = in_data[26079:26048] - in_data[26111:26080];
  assign out_data[130559:130528] = in_data[261087:261056] - in_data[261119:261088];
  assign out_data[130591:130560] = in_data[261151:261120] - in_data[261183:261152];
  assign out_data[130623:130592] = in_data[261215:261184] - in_data[261247:261216];
  assign out_data[130655:130624] = in_data[261279:261248] - in_data[261311:261280];
  assign out_data[130687:130656] = in_data[261343:261312] - in_data[261375:261344];
  assign out_data[130719:130688] = in_data[261407:261376] - in_data[261439:261408];
  assign out_data[130751:130720] = in_data[261471:261440] - in_data[261503:261472];
  assign out_data[130783:130752] = in_data[261535:261504] - in_data[261567:261536];
  assign out_data[130815:130784] = in_data[261599:261568] - in_data[261631:261600];
  assign out_data[130847:130816] = in_data[261663:261632] - in_data[261695:261664];
  assign out_data[13087:13056] = in_data[26143:26112] - in_data[26175:26144];
  assign out_data[130879:130848] = in_data[261727:261696] - in_data[261759:261728];
  assign out_data[130911:130880] = in_data[261791:261760] - in_data[261823:261792];
  assign out_data[130943:130912] = in_data[261855:261824] - in_data[261887:261856];
  assign out_data[130975:130944] = in_data[261919:261888] - in_data[261951:261920];
  assign out_data[131007:130976] = in_data[261983:261952] - in_data[262015:261984];
  assign out_data[131039:131008] = in_data[262047:262016] - in_data[262079:262048];
  assign out_data[131071:131040] = in_data[262111:262080] - in_data[262143:262112];
  assign out_data[1311:1280] = in_data[2591:2560] - in_data[2623:2592];
  assign out_data[13119:13088] = in_data[26207:26176] - in_data[26239:26208];
  assign out_data[13151:13120] = in_data[26271:26240] - in_data[26303:26272];
  assign out_data[13183:13152] = in_data[26335:26304] - in_data[26367:26336];
  assign out_data[13215:13184] = in_data[26399:26368] - in_data[26431:26400];
  assign out_data[13247:13216] = in_data[26463:26432] - in_data[26495:26464];
  assign out_data[13279:13248] = in_data[26527:26496] - in_data[26559:26528];
  assign out_data[13311:13280] = in_data[26591:26560] - in_data[26623:26592];
  assign out_data[13343:13312] = in_data[26655:26624] - in_data[26687:26656];
  assign out_data[13375:13344] = in_data[26719:26688] - in_data[26751:26720];
  assign out_data[13407:13376] = in_data[26783:26752] - in_data[26815:26784];
  assign out_data[1343:1312] = in_data[2655:2624] - in_data[2687:2656];
  assign out_data[13439:13408] = in_data[26847:26816] - in_data[26879:26848];
  assign out_data[13471:13440] = in_data[26911:26880] - in_data[26943:26912];
  assign out_data[13503:13472] = in_data[26975:26944] - in_data[27007:26976];
  assign out_data[13535:13504] = in_data[27039:27008] - in_data[27071:27040];
  assign out_data[13567:13536] = in_data[27103:27072] - in_data[27135:27104];
  assign out_data[13599:13568] = in_data[27167:27136] - in_data[27199:27168];
  assign out_data[13631:13600] = in_data[27231:27200] - in_data[27263:27232];
  assign out_data[13663:13632] = in_data[27295:27264] - in_data[27327:27296];
  assign out_data[13695:13664] = in_data[27359:27328] - in_data[27391:27360];
  assign out_data[13727:13696] = in_data[27423:27392] - in_data[27455:27424];
  assign out_data[1375:1344] = in_data[2719:2688] - in_data[2751:2720];
  assign out_data[13759:13728] = in_data[27487:27456] - in_data[27519:27488];
  assign out_data[13791:13760] = in_data[27551:27520] - in_data[27583:27552];
  assign out_data[13823:13792] = in_data[27615:27584] - in_data[27647:27616];
  assign out_data[13855:13824] = in_data[27679:27648] - in_data[27711:27680];
  assign out_data[13887:13856] = in_data[27743:27712] - in_data[27775:27744];
  assign out_data[13919:13888] = in_data[27807:27776] - in_data[27839:27808];
  assign out_data[13951:13920] = in_data[27871:27840] - in_data[27903:27872];
  assign out_data[13983:13952] = in_data[27935:27904] - in_data[27967:27936];
  assign out_data[14015:13984] = in_data[27999:27968] - in_data[28031:28000];
  assign out_data[14047:14016] = in_data[28063:28032] - in_data[28095:28064];
  assign out_data[1407:1376] = in_data[2783:2752] - in_data[2815:2784];
  assign out_data[14079:14048] = in_data[28127:28096] - in_data[28159:28128];
  assign out_data[14111:14080] = in_data[28191:28160] - in_data[28223:28192];
  assign out_data[14143:14112] = in_data[28255:28224] - in_data[28287:28256];
  assign out_data[14175:14144] = in_data[28319:28288] - in_data[28351:28320];
  assign out_data[14207:14176] = in_data[28383:28352] - in_data[28415:28384];
  assign out_data[14239:14208] = in_data[28447:28416] - in_data[28479:28448];
  assign out_data[14271:14240] = in_data[28511:28480] - in_data[28543:28512];
  assign out_data[14303:14272] = in_data[28575:28544] - in_data[28607:28576];
  assign out_data[14335:14304] = in_data[28639:28608] - in_data[28671:28640];
  assign out_data[14367:14336] = in_data[28703:28672] - in_data[28735:28704];
  assign out_data[1439:1408] = in_data[2847:2816] - in_data[2879:2848];
  assign out_data[14399:14368] = in_data[28767:28736] - in_data[28799:28768];
  assign out_data[14431:14400] = in_data[28831:28800] - in_data[28863:28832];
  assign out_data[14463:14432] = in_data[28895:28864] - in_data[28927:28896];
  assign out_data[14495:14464] = in_data[28959:28928] - in_data[28991:28960];
  assign out_data[14527:14496] = in_data[29023:28992] - in_data[29055:29024];
  assign out_data[14559:14528] = in_data[29087:29056] - in_data[29119:29088];
  assign out_data[14591:14560] = in_data[29151:29120] - in_data[29183:29152];
  assign out_data[14623:14592] = in_data[29215:29184] - in_data[29247:29216];
  assign out_data[14655:14624] = in_data[29279:29248] - in_data[29311:29280];
  assign out_data[14687:14656] = in_data[29343:29312] - in_data[29375:29344];
  assign out_data[1471:1440] = in_data[2911:2880] - in_data[2943:2912];
  assign out_data[14719:14688] = in_data[29407:29376] - in_data[29439:29408];
  assign out_data[14751:14720] = in_data[29471:29440] - in_data[29503:29472];
  assign out_data[14783:14752] = in_data[29535:29504] - in_data[29567:29536];
  assign out_data[14815:14784] = in_data[29599:29568] - in_data[29631:29600];
  assign out_data[14847:14816] = in_data[29663:29632] - in_data[29695:29664];
  assign out_data[14879:14848] = in_data[29727:29696] - in_data[29759:29728];
  assign out_data[14911:14880] = in_data[29791:29760] - in_data[29823:29792];
  assign out_data[14943:14912] = in_data[29855:29824] - in_data[29887:29856];
  assign out_data[14975:14944] = in_data[29919:29888] - in_data[29951:29920];
  assign out_data[15007:14976] = in_data[29983:29952] - in_data[30015:29984];
  assign out_data[1503:1472] = in_data[2975:2944] - in_data[3007:2976];
  assign out_data[15039:15008] = in_data[30047:30016] - in_data[30079:30048];
  assign out_data[15071:15040] = in_data[30111:30080] - in_data[30143:30112];
  assign out_data[15103:15072] = in_data[30175:30144] - in_data[30207:30176];
  assign out_data[15135:15104] = in_data[30239:30208] - in_data[30271:30240];
  assign out_data[15167:15136] = in_data[30303:30272] - in_data[30335:30304];
  assign out_data[15199:15168] = in_data[30367:30336] - in_data[30399:30368];
  assign out_data[15231:15200] = in_data[30431:30400] - in_data[30463:30432];
  assign out_data[15263:15232] = in_data[30495:30464] - in_data[30527:30496];
  assign out_data[15295:15264] = in_data[30559:30528] - in_data[30591:30560];
  assign out_data[15327:15296] = in_data[30623:30592] - in_data[30655:30624];
  assign out_data[1535:1504] = in_data[3039:3008] - in_data[3071:3040];
  assign out_data[15359:15328] = in_data[30687:30656] - in_data[30719:30688];
  assign out_data[15391:15360] = in_data[30751:30720] - in_data[30783:30752];
  assign out_data[15423:15392] = in_data[30815:30784] - in_data[30847:30816];
  assign out_data[15455:15424] = in_data[30879:30848] - in_data[30911:30880];
  assign out_data[15487:15456] = in_data[30943:30912] - in_data[30975:30944];
  assign out_data[15519:15488] = in_data[31007:30976] - in_data[31039:31008];
  assign out_data[15551:15520] = in_data[31071:31040] - in_data[31103:31072];
  assign out_data[15583:15552] = in_data[31135:31104] - in_data[31167:31136];
  assign out_data[15615:15584] = in_data[31199:31168] - in_data[31231:31200];
  assign out_data[15647:15616] = in_data[31263:31232] - in_data[31295:31264];
  assign out_data[1567:1536] = in_data[3103:3072] - in_data[3135:3104];
  assign out_data[15679:15648] = in_data[31327:31296] - in_data[31359:31328];
  assign out_data[15711:15680] = in_data[31391:31360] - in_data[31423:31392];
  assign out_data[15743:15712] = in_data[31455:31424] - in_data[31487:31456];
  assign out_data[15775:15744] = in_data[31519:31488] - in_data[31551:31520];
  assign out_data[15807:15776] = in_data[31583:31552] - in_data[31615:31584];
  assign out_data[15839:15808] = in_data[31647:31616] - in_data[31679:31648];
  assign out_data[15871:15840] = in_data[31711:31680] - in_data[31743:31712];
  assign out_data[15903:15872] = in_data[31775:31744] - in_data[31807:31776];
  assign out_data[15935:15904] = in_data[31839:31808] - in_data[31871:31840];
  assign out_data[15967:15936] = in_data[31903:31872] - in_data[31935:31904];
  assign out_data[159:128] = in_data[287:256] - in_data[319:288];
  assign out_data[1599:1568] = in_data[3167:3136] - in_data[3199:3168];
  assign out_data[15999:15968] = in_data[31967:31936] - in_data[31999:31968];
  assign out_data[16031:16000] = in_data[32031:32000] - in_data[32063:32032];
  assign out_data[16063:16032] = in_data[32095:32064] - in_data[32127:32096];
  assign out_data[16095:16064] = in_data[32159:32128] - in_data[32191:32160];
  assign out_data[16127:16096] = in_data[32223:32192] - in_data[32255:32224];
  assign out_data[16159:16128] = in_data[32287:32256] - in_data[32319:32288];
  assign out_data[16191:16160] = in_data[32351:32320] - in_data[32383:32352];
  assign out_data[16223:16192] = in_data[32415:32384] - in_data[32447:32416];
  assign out_data[16255:16224] = in_data[32479:32448] - in_data[32511:32480];
  assign out_data[16287:16256] = in_data[32543:32512] - in_data[32575:32544];
  assign out_data[1631:1600] = in_data[3231:3200] - in_data[3263:3232];
  assign out_data[16319:16288] = in_data[32607:32576] - in_data[32639:32608];
  assign out_data[16351:16320] = in_data[32671:32640] - in_data[32703:32672];
  assign out_data[16383:16352] = in_data[32735:32704] - in_data[32767:32736];
  assign out_data[16415:16384] = in_data[32799:32768] - in_data[32831:32800];
  assign out_data[16447:16416] = in_data[32863:32832] - in_data[32895:32864];
  assign out_data[16479:16448] = in_data[32927:32896] - in_data[32959:32928];
  assign out_data[16511:16480] = in_data[32991:32960] - in_data[33023:32992];
  assign out_data[16543:16512] = in_data[33055:33024] - in_data[33087:33056];
  assign out_data[16575:16544] = in_data[33119:33088] - in_data[33151:33120];
  assign out_data[16607:16576] = in_data[33183:33152] - in_data[33215:33184];
  assign out_data[1663:1632] = in_data[3295:3264] - in_data[3327:3296];
  assign out_data[16639:16608] = in_data[33247:33216] - in_data[33279:33248];
  assign out_data[16671:16640] = in_data[33311:33280] - in_data[33343:33312];
  assign out_data[16703:16672] = in_data[33375:33344] - in_data[33407:33376];
  assign out_data[16735:16704] = in_data[33439:33408] - in_data[33471:33440];
  assign out_data[16767:16736] = in_data[33503:33472] - in_data[33535:33504];
  assign out_data[16799:16768] = in_data[33567:33536] - in_data[33599:33568];
  assign out_data[16831:16800] = in_data[33631:33600] - in_data[33663:33632];
  assign out_data[16863:16832] = in_data[33695:33664] - in_data[33727:33696];
  assign out_data[16895:16864] = in_data[33759:33728] - in_data[33791:33760];
  assign out_data[16927:16896] = in_data[33823:33792] - in_data[33855:33824];
  assign out_data[1695:1664] = in_data[3359:3328] - in_data[3391:3360];
  assign out_data[16959:16928] = in_data[33887:33856] - in_data[33919:33888];
  assign out_data[16991:16960] = in_data[33951:33920] - in_data[33983:33952];
  assign out_data[17023:16992] = in_data[34015:33984] - in_data[34047:34016];
  assign out_data[17055:17024] = in_data[34079:34048] - in_data[34111:34080];
  assign out_data[17087:17056] = in_data[34143:34112] - in_data[34175:34144];
  assign out_data[17119:17088] = in_data[34207:34176] - in_data[34239:34208];
  assign out_data[17151:17120] = in_data[34271:34240] - in_data[34303:34272];
  assign out_data[17183:17152] = in_data[34335:34304] - in_data[34367:34336];
  assign out_data[17215:17184] = in_data[34399:34368] - in_data[34431:34400];
  assign out_data[17247:17216] = in_data[34463:34432] - in_data[34495:34464];
  assign out_data[1727:1696] = in_data[3423:3392] - in_data[3455:3424];
  assign out_data[17279:17248] = in_data[34527:34496] - in_data[34559:34528];
  assign out_data[17311:17280] = in_data[34591:34560] - in_data[34623:34592];
  assign out_data[17343:17312] = in_data[34655:34624] - in_data[34687:34656];
  assign out_data[17375:17344] = in_data[34719:34688] - in_data[34751:34720];
  assign out_data[17407:17376] = in_data[34783:34752] - in_data[34815:34784];
  assign out_data[17439:17408] = in_data[34847:34816] - in_data[34879:34848];
  assign out_data[17471:17440] = in_data[34911:34880] - in_data[34943:34912];
  assign out_data[17503:17472] = in_data[34975:34944] - in_data[35007:34976];
  assign out_data[17535:17504] = in_data[35039:35008] - in_data[35071:35040];
  assign out_data[17567:17536] = in_data[35103:35072] - in_data[35135:35104];
  assign out_data[1759:1728] = in_data[3487:3456] - in_data[3519:3488];
  assign out_data[17599:17568] = in_data[35167:35136] - in_data[35199:35168];
  assign out_data[17631:17600] = in_data[35231:35200] - in_data[35263:35232];
  assign out_data[17663:17632] = in_data[35295:35264] - in_data[35327:35296];
  assign out_data[17695:17664] = in_data[35359:35328] - in_data[35391:35360];
  assign out_data[17727:17696] = in_data[35423:35392] - in_data[35455:35424];
  assign out_data[17759:17728] = in_data[35487:35456] - in_data[35519:35488];
  assign out_data[17791:17760] = in_data[35551:35520] - in_data[35583:35552];
  assign out_data[17823:17792] = in_data[35615:35584] - in_data[35647:35616];
  assign out_data[17855:17824] = in_data[35679:35648] - in_data[35711:35680];
  assign out_data[17887:17856] = in_data[35743:35712] - in_data[35775:35744];
  assign out_data[1791:1760] = in_data[3551:3520] - in_data[3583:3552];
  assign out_data[17919:17888] = in_data[35807:35776] - in_data[35839:35808];
  assign out_data[17951:17920] = in_data[35871:35840] - in_data[35903:35872];
  assign out_data[17983:17952] = in_data[35935:35904] - in_data[35967:35936];
  assign out_data[18015:17984] = in_data[35999:35968] - in_data[36031:36000];
  assign out_data[18047:18016] = in_data[36063:36032] - in_data[36095:36064];
  assign out_data[18079:18048] = in_data[36127:36096] - in_data[36159:36128];
  assign out_data[18111:18080] = in_data[36191:36160] - in_data[36223:36192];
  assign out_data[18143:18112] = in_data[36255:36224] - in_data[36287:36256];
  assign out_data[18175:18144] = in_data[36319:36288] - in_data[36351:36320];
  assign out_data[18207:18176] = in_data[36383:36352] - in_data[36415:36384];
  assign out_data[1823:1792] = in_data[3615:3584] - in_data[3647:3616];
  assign out_data[18239:18208] = in_data[36447:36416] - in_data[36479:36448];
  assign out_data[18271:18240] = in_data[36511:36480] - in_data[36543:36512];
  assign out_data[18303:18272] = in_data[36575:36544] - in_data[36607:36576];
  assign out_data[18335:18304] = in_data[36639:36608] - in_data[36671:36640];
  assign out_data[18367:18336] = in_data[36703:36672] - in_data[36735:36704];
  assign out_data[18399:18368] = in_data[36767:36736] - in_data[36799:36768];
  assign out_data[18431:18400] = in_data[36831:36800] - in_data[36863:36832];
  assign out_data[18463:18432] = in_data[36895:36864] - in_data[36927:36896];
  assign out_data[18495:18464] = in_data[36959:36928] - in_data[36991:36960];
  assign out_data[18527:18496] = in_data[37023:36992] - in_data[37055:37024];
  assign out_data[1855:1824] = in_data[3679:3648] - in_data[3711:3680];
  assign out_data[18559:18528] = in_data[37087:37056] - in_data[37119:37088];
  assign out_data[18591:18560] = in_data[37151:37120] - in_data[37183:37152];
  assign out_data[18623:18592] = in_data[37215:37184] - in_data[37247:37216];
  assign out_data[18655:18624] = in_data[37279:37248] - in_data[37311:37280];
  assign out_data[18687:18656] = in_data[37343:37312] - in_data[37375:37344];
  assign out_data[18719:18688] = in_data[37407:37376] - in_data[37439:37408];
  assign out_data[18751:18720] = in_data[37471:37440] - in_data[37503:37472];
  assign out_data[18783:18752] = in_data[37535:37504] - in_data[37567:37536];
  assign out_data[18815:18784] = in_data[37599:37568] - in_data[37631:37600];
  assign out_data[18847:18816] = in_data[37663:37632] - in_data[37695:37664];
  assign out_data[1887:1856] = in_data[3743:3712] - in_data[3775:3744];
  assign out_data[18879:18848] = in_data[37727:37696] - in_data[37759:37728];
  assign out_data[18911:18880] = in_data[37791:37760] - in_data[37823:37792];
  assign out_data[18943:18912] = in_data[37855:37824] - in_data[37887:37856];
  assign out_data[18975:18944] = in_data[37919:37888] - in_data[37951:37920];
  assign out_data[19007:18976] = in_data[37983:37952] - in_data[38015:37984];
  assign out_data[19039:19008] = in_data[38047:38016] - in_data[38079:38048];
  assign out_data[19071:19040] = in_data[38111:38080] - in_data[38143:38112];
  assign out_data[19103:19072] = in_data[38175:38144] - in_data[38207:38176];
  assign out_data[19135:19104] = in_data[38239:38208] - in_data[38271:38240];
  assign out_data[19167:19136] = in_data[38303:38272] - in_data[38335:38304];
  assign out_data[191:160] = in_data[351:320] - in_data[383:352];
  assign out_data[1919:1888] = in_data[3807:3776] - in_data[3839:3808];
  assign out_data[19199:19168] = in_data[38367:38336] - in_data[38399:38368];
  assign out_data[19231:19200] = in_data[38431:38400] - in_data[38463:38432];
  assign out_data[19263:19232] = in_data[38495:38464] - in_data[38527:38496];
  assign out_data[19295:19264] = in_data[38559:38528] - in_data[38591:38560];
  assign out_data[19327:19296] = in_data[38623:38592] - in_data[38655:38624];
  assign out_data[19359:19328] = in_data[38687:38656] - in_data[38719:38688];
  assign out_data[19391:19360] = in_data[38751:38720] - in_data[38783:38752];
  assign out_data[19423:19392] = in_data[38815:38784] - in_data[38847:38816];
  assign out_data[19455:19424] = in_data[38879:38848] - in_data[38911:38880];
  assign out_data[19487:19456] = in_data[38943:38912] - in_data[38975:38944];
  assign out_data[1951:1920] = in_data[3871:3840] - in_data[3903:3872];
  assign out_data[19519:19488] = in_data[39007:38976] - in_data[39039:39008];
  assign out_data[19551:19520] = in_data[39071:39040] - in_data[39103:39072];
  assign out_data[19583:19552] = in_data[39135:39104] - in_data[39167:39136];
  assign out_data[19615:19584] = in_data[39199:39168] - in_data[39231:39200];
  assign out_data[19647:19616] = in_data[39263:39232] - in_data[39295:39264];
  assign out_data[19679:19648] = in_data[39327:39296] - in_data[39359:39328];
  assign out_data[19711:19680] = in_data[39391:39360] - in_data[39423:39392];
  assign out_data[19743:19712] = in_data[39455:39424] - in_data[39487:39456];
  assign out_data[19775:19744] = in_data[39519:39488] - in_data[39551:39520];
  assign out_data[19807:19776] = in_data[39583:39552] - in_data[39615:39584];
  assign out_data[1983:1952] = in_data[3935:3904] - in_data[3967:3936];
  assign out_data[19839:19808] = in_data[39647:39616] - in_data[39679:39648];
  assign out_data[19871:19840] = in_data[39711:39680] - in_data[39743:39712];
  assign out_data[19903:19872] = in_data[39775:39744] - in_data[39807:39776];
  assign out_data[19935:19904] = in_data[39839:39808] - in_data[39871:39840];
  assign out_data[19967:19936] = in_data[39903:39872] - in_data[39935:39904];
  assign out_data[19999:19968] = in_data[39967:39936] - in_data[39999:39968];
  assign out_data[20031:20000] = in_data[40031:40000] - in_data[40063:40032];
  assign out_data[20063:20032] = in_data[40095:40064] - in_data[40127:40096];
  assign out_data[20095:20064] = in_data[40159:40128] - in_data[40191:40160];
  assign out_data[20127:20096] = in_data[40223:40192] - in_data[40255:40224];
  assign out_data[2015:1984] = in_data[3999:3968] - in_data[4031:4000];
  assign out_data[20159:20128] = in_data[40287:40256] - in_data[40319:40288];
  assign out_data[20191:20160] = in_data[40351:40320] - in_data[40383:40352];
  assign out_data[20223:20192] = in_data[40415:40384] - in_data[40447:40416];
  assign out_data[20255:20224] = in_data[40479:40448] - in_data[40511:40480];
  assign out_data[20287:20256] = in_data[40543:40512] - in_data[40575:40544];
  assign out_data[20319:20288] = in_data[40607:40576] - in_data[40639:40608];
  assign out_data[20351:20320] = in_data[40671:40640] - in_data[40703:40672];
  assign out_data[20383:20352] = in_data[40735:40704] - in_data[40767:40736];
  assign out_data[20415:20384] = in_data[40799:40768] - in_data[40831:40800];
  assign out_data[20447:20416] = in_data[40863:40832] - in_data[40895:40864];
  assign out_data[2047:2016] = in_data[4063:4032] - in_data[4095:4064];
  assign out_data[20479:20448] = in_data[40927:40896] - in_data[40959:40928];
  assign out_data[20511:20480] = in_data[40991:40960] - in_data[41023:40992];
  assign out_data[20543:20512] = in_data[41055:41024] - in_data[41087:41056];
  assign out_data[20575:20544] = in_data[41119:41088] - in_data[41151:41120];
  assign out_data[20607:20576] = in_data[41183:41152] - in_data[41215:41184];
  assign out_data[20639:20608] = in_data[41247:41216] - in_data[41279:41248];
  assign out_data[20671:20640] = in_data[41311:41280] - in_data[41343:41312];
  assign out_data[20703:20672] = in_data[41375:41344] - in_data[41407:41376];
  assign out_data[20735:20704] = in_data[41439:41408] - in_data[41471:41440];
  assign out_data[20767:20736] = in_data[41503:41472] - in_data[41535:41504];
  assign out_data[2079:2048] = in_data[4127:4096] - in_data[4159:4128];
  assign out_data[20799:20768] = in_data[41567:41536] - in_data[41599:41568];
  assign out_data[20831:20800] = in_data[41631:41600] - in_data[41663:41632];
  assign out_data[20863:20832] = in_data[41695:41664] - in_data[41727:41696];
  assign out_data[20895:20864] = in_data[41759:41728] - in_data[41791:41760];
  assign out_data[20927:20896] = in_data[41823:41792] - in_data[41855:41824];
  assign out_data[20959:20928] = in_data[41887:41856] - in_data[41919:41888];
  assign out_data[20991:20960] = in_data[41951:41920] - in_data[41983:41952];
  assign out_data[21023:20992] = in_data[42015:41984] - in_data[42047:42016];
  assign out_data[21055:21024] = in_data[42079:42048] - in_data[42111:42080];
  assign out_data[21087:21056] = in_data[42143:42112] - in_data[42175:42144];
  assign out_data[2111:2080] = in_data[4191:4160] - in_data[4223:4192];
  assign out_data[21119:21088] = in_data[42207:42176] - in_data[42239:42208];
  assign out_data[21151:21120] = in_data[42271:42240] - in_data[42303:42272];
  assign out_data[21183:21152] = in_data[42335:42304] - in_data[42367:42336];
  assign out_data[21215:21184] = in_data[42399:42368] - in_data[42431:42400];
  assign out_data[21247:21216] = in_data[42463:42432] - in_data[42495:42464];
  assign out_data[21279:21248] = in_data[42527:42496] - in_data[42559:42528];
  assign out_data[21311:21280] = in_data[42591:42560] - in_data[42623:42592];
  assign out_data[21343:21312] = in_data[42655:42624] - in_data[42687:42656];
  assign out_data[21375:21344] = in_data[42719:42688] - in_data[42751:42720];
  assign out_data[21407:21376] = in_data[42783:42752] - in_data[42815:42784];
  assign out_data[2143:2112] = in_data[4255:4224] - in_data[4287:4256];
  assign out_data[21439:21408] = in_data[42847:42816] - in_data[42879:42848];
  assign out_data[21471:21440] = in_data[42911:42880] - in_data[42943:42912];
  assign out_data[21503:21472] = in_data[42975:42944] - in_data[43007:42976];
  assign out_data[21535:21504] = in_data[43039:43008] - in_data[43071:43040];
  assign out_data[21567:21536] = in_data[43103:43072] - in_data[43135:43104];
  assign out_data[21599:21568] = in_data[43167:43136] - in_data[43199:43168];
  assign out_data[21631:21600] = in_data[43231:43200] - in_data[43263:43232];
  assign out_data[21663:21632] = in_data[43295:43264] - in_data[43327:43296];
  assign out_data[21695:21664] = in_data[43359:43328] - in_data[43391:43360];
  assign out_data[21727:21696] = in_data[43423:43392] - in_data[43455:43424];
  assign out_data[2175:2144] = in_data[4319:4288] - in_data[4351:4320];
  assign out_data[21759:21728] = in_data[43487:43456] - in_data[43519:43488];
  assign out_data[21791:21760] = in_data[43551:43520] - in_data[43583:43552];
  assign out_data[21823:21792] = in_data[43615:43584] - in_data[43647:43616];
  assign out_data[21855:21824] = in_data[43679:43648] - in_data[43711:43680];
  assign out_data[21887:21856] = in_data[43743:43712] - in_data[43775:43744];
  assign out_data[21919:21888] = in_data[43807:43776] - in_data[43839:43808];
  assign out_data[21951:21920] = in_data[43871:43840] - in_data[43903:43872];
  assign out_data[21983:21952] = in_data[43935:43904] - in_data[43967:43936];
  assign out_data[22015:21984] = in_data[43999:43968] - in_data[44031:44000];
  assign out_data[22047:22016] = in_data[44063:44032] - in_data[44095:44064];
  assign out_data[2207:2176] = in_data[4383:4352] - in_data[4415:4384];
  assign out_data[22079:22048] = in_data[44127:44096] - in_data[44159:44128];
  assign out_data[22111:22080] = in_data[44191:44160] - in_data[44223:44192];
  assign out_data[22143:22112] = in_data[44255:44224] - in_data[44287:44256];
  assign out_data[22175:22144] = in_data[44319:44288] - in_data[44351:44320];
  assign out_data[22207:22176] = in_data[44383:44352] - in_data[44415:44384];
  assign out_data[22239:22208] = in_data[44447:44416] - in_data[44479:44448];
  assign out_data[22271:22240] = in_data[44511:44480] - in_data[44543:44512];
  assign out_data[22303:22272] = in_data[44575:44544] - in_data[44607:44576];
  assign out_data[22335:22304] = in_data[44639:44608] - in_data[44671:44640];
  assign out_data[22367:22336] = in_data[44703:44672] - in_data[44735:44704];
  assign out_data[223:192] = in_data[415:384] - in_data[447:416];
  assign out_data[2239:2208] = in_data[4447:4416] - in_data[4479:4448];
  assign out_data[22399:22368] = in_data[44767:44736] - in_data[44799:44768];
  assign out_data[22431:22400] = in_data[44831:44800] - in_data[44863:44832];
  assign out_data[22463:22432] = in_data[44895:44864] - in_data[44927:44896];
  assign out_data[22495:22464] = in_data[44959:44928] - in_data[44991:44960];
  assign out_data[22527:22496] = in_data[45023:44992] - in_data[45055:45024];
  assign out_data[22559:22528] = in_data[45087:45056] - in_data[45119:45088];
  assign out_data[22591:22560] = in_data[45151:45120] - in_data[45183:45152];
  assign out_data[22623:22592] = in_data[45215:45184] - in_data[45247:45216];
  assign out_data[22655:22624] = in_data[45279:45248] - in_data[45311:45280];
  assign out_data[22687:22656] = in_data[45343:45312] - in_data[45375:45344];
  assign out_data[2271:2240] = in_data[4511:4480] - in_data[4543:4512];
  assign out_data[22719:22688] = in_data[45407:45376] - in_data[45439:45408];
  assign out_data[22751:22720] = in_data[45471:45440] - in_data[45503:45472];
  assign out_data[22783:22752] = in_data[45535:45504] - in_data[45567:45536];
  assign out_data[22815:22784] = in_data[45599:45568] - in_data[45631:45600];
  assign out_data[22847:22816] = in_data[45663:45632] - in_data[45695:45664];
  assign out_data[22879:22848] = in_data[45727:45696] - in_data[45759:45728];
  assign out_data[22911:22880] = in_data[45791:45760] - in_data[45823:45792];
  assign out_data[22943:22912] = in_data[45855:45824] - in_data[45887:45856];
  assign out_data[22975:22944] = in_data[45919:45888] - in_data[45951:45920];
  assign out_data[23007:22976] = in_data[45983:45952] - in_data[46015:45984];
  assign out_data[2303:2272] = in_data[4575:4544] - in_data[4607:4576];
  assign out_data[23039:23008] = in_data[46047:46016] - in_data[46079:46048];
  assign out_data[23071:23040] = in_data[46111:46080] - in_data[46143:46112];
  assign out_data[23103:23072] = in_data[46175:46144] - in_data[46207:46176];
  assign out_data[23135:23104] = in_data[46239:46208] - in_data[46271:46240];
  assign out_data[23167:23136] = in_data[46303:46272] - in_data[46335:46304];
  assign out_data[23199:23168] = in_data[46367:46336] - in_data[46399:46368];
  assign out_data[23231:23200] = in_data[46431:46400] - in_data[46463:46432];
  assign out_data[23263:23232] = in_data[46495:46464] - in_data[46527:46496];
  assign out_data[23295:23264] = in_data[46559:46528] - in_data[46591:46560];
  assign out_data[23327:23296] = in_data[46623:46592] - in_data[46655:46624];
  assign out_data[2335:2304] = in_data[4639:4608] - in_data[4671:4640];
  assign out_data[23359:23328] = in_data[46687:46656] - in_data[46719:46688];
  assign out_data[23391:23360] = in_data[46751:46720] - in_data[46783:46752];
  assign out_data[23423:23392] = in_data[46815:46784] - in_data[46847:46816];
  assign out_data[23455:23424] = in_data[46879:46848] - in_data[46911:46880];
  assign out_data[23487:23456] = in_data[46943:46912] - in_data[46975:46944];
  assign out_data[23519:23488] = in_data[47007:46976] - in_data[47039:47008];
  assign out_data[23551:23520] = in_data[47071:47040] - in_data[47103:47072];
  assign out_data[23583:23552] = in_data[47135:47104] - in_data[47167:47136];
  assign out_data[23615:23584] = in_data[47199:47168] - in_data[47231:47200];
  assign out_data[23647:23616] = in_data[47263:47232] - in_data[47295:47264];
  assign out_data[2367:2336] = in_data[4703:4672] - in_data[4735:4704];
  assign out_data[23679:23648] = in_data[47327:47296] - in_data[47359:47328];
  assign out_data[23711:23680] = in_data[47391:47360] - in_data[47423:47392];
  assign out_data[23743:23712] = in_data[47455:47424] - in_data[47487:47456];
  assign out_data[23775:23744] = in_data[47519:47488] - in_data[47551:47520];
  assign out_data[23807:23776] = in_data[47583:47552] - in_data[47615:47584];
  assign out_data[23839:23808] = in_data[47647:47616] - in_data[47679:47648];
  assign out_data[23871:23840] = in_data[47711:47680] - in_data[47743:47712];
  assign out_data[23903:23872] = in_data[47775:47744] - in_data[47807:47776];
  assign out_data[23935:23904] = in_data[47839:47808] - in_data[47871:47840];
  assign out_data[23967:23936] = in_data[47903:47872] - in_data[47935:47904];
  assign out_data[2399:2368] = in_data[4767:4736] - in_data[4799:4768];
  assign out_data[23999:23968] = in_data[47967:47936] - in_data[47999:47968];
  assign out_data[24031:24000] = in_data[48031:48000] - in_data[48063:48032];
  assign out_data[24063:24032] = in_data[48095:48064] - in_data[48127:48096];
  assign out_data[24095:24064] = in_data[48159:48128] - in_data[48191:48160];
  assign out_data[24127:24096] = in_data[48223:48192] - in_data[48255:48224];
  assign out_data[24159:24128] = in_data[48287:48256] - in_data[48319:48288];
  assign out_data[24191:24160] = in_data[48351:48320] - in_data[48383:48352];
  assign out_data[24223:24192] = in_data[48415:48384] - in_data[48447:48416];
  assign out_data[24255:24224] = in_data[48479:48448] - in_data[48511:48480];
  assign out_data[24287:24256] = in_data[48543:48512] - in_data[48575:48544];
  assign out_data[2431:2400] = in_data[4831:4800] - in_data[4863:4832];
  assign out_data[24319:24288] = in_data[48607:48576] - in_data[48639:48608];
  assign out_data[24351:24320] = in_data[48671:48640] - in_data[48703:48672];
  assign out_data[24383:24352] = in_data[48735:48704] - in_data[48767:48736];
  assign out_data[24415:24384] = in_data[48799:48768] - in_data[48831:48800];
  assign out_data[24447:24416] = in_data[48863:48832] - in_data[48895:48864];
  assign out_data[24479:24448] = in_data[48927:48896] - in_data[48959:48928];
  assign out_data[24511:24480] = in_data[48991:48960] - in_data[49023:48992];
  assign out_data[24543:24512] = in_data[49055:49024] - in_data[49087:49056];
  assign out_data[24575:24544] = in_data[49119:49088] - in_data[49151:49120];
  assign out_data[24607:24576] = in_data[49183:49152] - in_data[49215:49184];
  assign out_data[2463:2432] = in_data[4895:4864] - in_data[4927:4896];
  assign out_data[24639:24608] = in_data[49247:49216] - in_data[49279:49248];
  assign out_data[24671:24640] = in_data[49311:49280] - in_data[49343:49312];
  assign out_data[24703:24672] = in_data[49375:49344] - in_data[49407:49376];
  assign out_data[24735:24704] = in_data[49439:49408] - in_data[49471:49440];
  assign out_data[24767:24736] = in_data[49503:49472] - in_data[49535:49504];
  assign out_data[24799:24768] = in_data[49567:49536] - in_data[49599:49568];
  assign out_data[24831:24800] = in_data[49631:49600] - in_data[49663:49632];
  assign out_data[24863:24832] = in_data[49695:49664] - in_data[49727:49696];
  assign out_data[24895:24864] = in_data[49759:49728] - in_data[49791:49760];
  assign out_data[24927:24896] = in_data[49823:49792] - in_data[49855:49824];
  assign out_data[2495:2464] = in_data[4959:4928] - in_data[4991:4960];
  assign out_data[24959:24928] = in_data[49887:49856] - in_data[49919:49888];
  assign out_data[24991:24960] = in_data[49951:49920] - in_data[49983:49952];
  assign out_data[25023:24992] = in_data[50015:49984] - in_data[50047:50016];
  assign out_data[25055:25024] = in_data[50079:50048] - in_data[50111:50080];
  assign out_data[25087:25056] = in_data[50143:50112] - in_data[50175:50144];
  assign out_data[25119:25088] = in_data[50207:50176] - in_data[50239:50208];
  assign out_data[25151:25120] = in_data[50271:50240] - in_data[50303:50272];
  assign out_data[25183:25152] = in_data[50335:50304] - in_data[50367:50336];
  assign out_data[25215:25184] = in_data[50399:50368] - in_data[50431:50400];
  assign out_data[25247:25216] = in_data[50463:50432] - in_data[50495:50464];
  assign out_data[2527:2496] = in_data[5023:4992] - in_data[5055:5024];
  assign out_data[25279:25248] = in_data[50527:50496] - in_data[50559:50528];
  assign out_data[25311:25280] = in_data[50591:50560] - in_data[50623:50592];
  assign out_data[25343:25312] = in_data[50655:50624] - in_data[50687:50656];
  assign out_data[25375:25344] = in_data[50719:50688] - in_data[50751:50720];
  assign out_data[25407:25376] = in_data[50783:50752] - in_data[50815:50784];
  assign out_data[25439:25408] = in_data[50847:50816] - in_data[50879:50848];
  assign out_data[25471:25440] = in_data[50911:50880] - in_data[50943:50912];
  assign out_data[25503:25472] = in_data[50975:50944] - in_data[51007:50976];
  assign out_data[25535:25504] = in_data[51039:51008] - in_data[51071:51040];
  assign out_data[25567:25536] = in_data[51103:51072] - in_data[51135:51104];
  assign out_data[255:224] = in_data[479:448] - in_data[511:480];
  assign out_data[2559:2528] = in_data[5087:5056] - in_data[5119:5088];
  assign out_data[25599:25568] = in_data[51167:51136] - in_data[51199:51168];
  assign out_data[25631:25600] = in_data[51231:51200] - in_data[51263:51232];
  assign out_data[25663:25632] = in_data[51295:51264] - in_data[51327:51296];
  assign out_data[25695:25664] = in_data[51359:51328] - in_data[51391:51360];
  assign out_data[25727:25696] = in_data[51423:51392] - in_data[51455:51424];
  assign out_data[25759:25728] = in_data[51487:51456] - in_data[51519:51488];
  assign out_data[25791:25760] = in_data[51551:51520] - in_data[51583:51552];
  assign out_data[25823:25792] = in_data[51615:51584] - in_data[51647:51616];
  assign out_data[25855:25824] = in_data[51679:51648] - in_data[51711:51680];
  assign out_data[25887:25856] = in_data[51743:51712] - in_data[51775:51744];
  assign out_data[2591:2560] = in_data[5151:5120] - in_data[5183:5152];
  assign out_data[25919:25888] = in_data[51807:51776] - in_data[51839:51808];
  assign out_data[25951:25920] = in_data[51871:51840] - in_data[51903:51872];
  assign out_data[25983:25952] = in_data[51935:51904] - in_data[51967:51936];
  assign out_data[26015:25984] = in_data[51999:51968] - in_data[52031:52000];
  assign out_data[26047:26016] = in_data[52063:52032] - in_data[52095:52064];
  assign out_data[26079:26048] = in_data[52127:52096] - in_data[52159:52128];
  assign out_data[26111:26080] = in_data[52191:52160] - in_data[52223:52192];
  assign out_data[26143:26112] = in_data[52255:52224] - in_data[52287:52256];
  assign out_data[26175:26144] = in_data[52319:52288] - in_data[52351:52320];
  assign out_data[26207:26176] = in_data[52383:52352] - in_data[52415:52384];
  assign out_data[2623:2592] = in_data[5215:5184] - in_data[5247:5216];
  assign out_data[26239:26208] = in_data[52447:52416] - in_data[52479:52448];
  assign out_data[26271:26240] = in_data[52511:52480] - in_data[52543:52512];
  assign out_data[26303:26272] = in_data[52575:52544] - in_data[52607:52576];
  assign out_data[26335:26304] = in_data[52639:52608] - in_data[52671:52640];
  assign out_data[26367:26336] = in_data[52703:52672] - in_data[52735:52704];
  assign out_data[26399:26368] = in_data[52767:52736] - in_data[52799:52768];
  assign out_data[26431:26400] = in_data[52831:52800] - in_data[52863:52832];
  assign out_data[26463:26432] = in_data[52895:52864] - in_data[52927:52896];
  assign out_data[26495:26464] = in_data[52959:52928] - in_data[52991:52960];
  assign out_data[26527:26496] = in_data[53023:52992] - in_data[53055:53024];
  assign out_data[2655:2624] = in_data[5279:5248] - in_data[5311:5280];
  assign out_data[26559:26528] = in_data[53087:53056] - in_data[53119:53088];
  assign out_data[26591:26560] = in_data[53151:53120] - in_data[53183:53152];
  assign out_data[26623:26592] = in_data[53215:53184] - in_data[53247:53216];
  assign out_data[26655:26624] = in_data[53279:53248] - in_data[53311:53280];
  assign out_data[26687:26656] = in_data[53343:53312] - in_data[53375:53344];
  assign out_data[26719:26688] = in_data[53407:53376] - in_data[53439:53408];
  assign out_data[26751:26720] = in_data[53471:53440] - in_data[53503:53472];
  assign out_data[26783:26752] = in_data[53535:53504] - in_data[53567:53536];
  assign out_data[26815:26784] = in_data[53599:53568] - in_data[53631:53600];
  assign out_data[26847:26816] = in_data[53663:53632] - in_data[53695:53664];
  assign out_data[2687:2656] = in_data[5343:5312] - in_data[5375:5344];
  assign out_data[26879:26848] = in_data[53727:53696] - in_data[53759:53728];
  assign out_data[26911:26880] = in_data[53791:53760] - in_data[53823:53792];
  assign out_data[26943:26912] = in_data[53855:53824] - in_data[53887:53856];
  assign out_data[26975:26944] = in_data[53919:53888] - in_data[53951:53920];
  assign out_data[27007:26976] = in_data[53983:53952] - in_data[54015:53984];
  assign out_data[27039:27008] = in_data[54047:54016] - in_data[54079:54048];
  assign out_data[27071:27040] = in_data[54111:54080] - in_data[54143:54112];
  assign out_data[27103:27072] = in_data[54175:54144] - in_data[54207:54176];
  assign out_data[27135:27104] = in_data[54239:54208] - in_data[54271:54240];
  assign out_data[27167:27136] = in_data[54303:54272] - in_data[54335:54304];
  assign out_data[2719:2688] = in_data[5407:5376] - in_data[5439:5408];
  assign out_data[27199:27168] = in_data[54367:54336] - in_data[54399:54368];
  assign out_data[27231:27200] = in_data[54431:54400] - in_data[54463:54432];
  assign out_data[27263:27232] = in_data[54495:54464] - in_data[54527:54496];
  assign out_data[27295:27264] = in_data[54559:54528] - in_data[54591:54560];
  assign out_data[27327:27296] = in_data[54623:54592] - in_data[54655:54624];
  assign out_data[27359:27328] = in_data[54687:54656] - in_data[54719:54688];
  assign out_data[27391:27360] = in_data[54751:54720] - in_data[54783:54752];
  assign out_data[27423:27392] = in_data[54815:54784] - in_data[54847:54816];
  assign out_data[27455:27424] = in_data[54879:54848] - in_data[54911:54880];
  assign out_data[27487:27456] = in_data[54943:54912] - in_data[54975:54944];
  assign out_data[2751:2720] = in_data[5471:5440] - in_data[5503:5472];
  assign out_data[27519:27488] = in_data[55007:54976] - in_data[55039:55008];
  assign out_data[27551:27520] = in_data[55071:55040] - in_data[55103:55072];
  assign out_data[27583:27552] = in_data[55135:55104] - in_data[55167:55136];
  assign out_data[27615:27584] = in_data[55199:55168] - in_data[55231:55200];
  assign out_data[27647:27616] = in_data[55263:55232] - in_data[55295:55264];
  assign out_data[27679:27648] = in_data[55327:55296] - in_data[55359:55328];
  assign out_data[27711:27680] = in_data[55391:55360] - in_data[55423:55392];
  assign out_data[27743:27712] = in_data[55455:55424] - in_data[55487:55456];
  assign out_data[27775:27744] = in_data[55519:55488] - in_data[55551:55520];
  assign out_data[27807:27776] = in_data[55583:55552] - in_data[55615:55584];
  assign out_data[2783:2752] = in_data[5535:5504] - in_data[5567:5536];
  assign out_data[27839:27808] = in_data[55647:55616] - in_data[55679:55648];
  assign out_data[27871:27840] = in_data[55711:55680] - in_data[55743:55712];
  assign out_data[27903:27872] = in_data[55775:55744] - in_data[55807:55776];
  assign out_data[27935:27904] = in_data[55839:55808] - in_data[55871:55840];
  assign out_data[27967:27936] = in_data[55903:55872] - in_data[55935:55904];
  assign out_data[27999:27968] = in_data[55967:55936] - in_data[55999:55968];
  assign out_data[28031:28000] = in_data[56031:56000] - in_data[56063:56032];
  assign out_data[28063:28032] = in_data[56095:56064] - in_data[56127:56096];
  assign out_data[28095:28064] = in_data[56159:56128] - in_data[56191:56160];
  assign out_data[28127:28096] = in_data[56223:56192] - in_data[56255:56224];
  assign out_data[2815:2784] = in_data[5599:5568] - in_data[5631:5600];
  assign out_data[28159:28128] = in_data[56287:56256] - in_data[56319:56288];
  assign out_data[28191:28160] = in_data[56351:56320] - in_data[56383:56352];
  assign out_data[28223:28192] = in_data[56415:56384] - in_data[56447:56416];
  assign out_data[28255:28224] = in_data[56479:56448] - in_data[56511:56480];
  assign out_data[28287:28256] = in_data[56543:56512] - in_data[56575:56544];
  assign out_data[28319:28288] = in_data[56607:56576] - in_data[56639:56608];
  assign out_data[28351:28320] = in_data[56671:56640] - in_data[56703:56672];
  assign out_data[28383:28352] = in_data[56735:56704] - in_data[56767:56736];
  assign out_data[28415:28384] = in_data[56799:56768] - in_data[56831:56800];
  assign out_data[28447:28416] = in_data[56863:56832] - in_data[56895:56864];
  assign out_data[2847:2816] = in_data[5663:5632] - in_data[5695:5664];
  assign out_data[28479:28448] = in_data[56927:56896] - in_data[56959:56928];
  assign out_data[28511:28480] = in_data[56991:56960] - in_data[57023:56992];
  assign out_data[28543:28512] = in_data[57055:57024] - in_data[57087:57056];
  assign out_data[28575:28544] = in_data[57119:57088] - in_data[57151:57120];
  assign out_data[28607:28576] = in_data[57183:57152] - in_data[57215:57184];
  assign out_data[28639:28608] = in_data[57247:57216] - in_data[57279:57248];
  assign out_data[28671:28640] = in_data[57311:57280] - in_data[57343:57312];
  assign out_data[28703:28672] = in_data[57375:57344] - in_data[57407:57376];
  assign out_data[28735:28704] = in_data[57439:57408] - in_data[57471:57440];
  assign out_data[28767:28736] = in_data[57503:57472] - in_data[57535:57504];
  assign out_data[287:256] = in_data[543:512] - in_data[575:544];
  assign out_data[2879:2848] = in_data[5727:5696] - in_data[5759:5728];
  assign out_data[28799:28768] = in_data[57567:57536] - in_data[57599:57568];
  assign out_data[28831:28800] = in_data[57631:57600] - in_data[57663:57632];
  assign out_data[28863:28832] = in_data[57695:57664] - in_data[57727:57696];
  assign out_data[28895:28864] = in_data[57759:57728] - in_data[57791:57760];
  assign out_data[28927:28896] = in_data[57823:57792] - in_data[57855:57824];
  assign out_data[28959:28928] = in_data[57887:57856] - in_data[57919:57888];
  assign out_data[28991:28960] = in_data[57951:57920] - in_data[57983:57952];
  assign out_data[29023:28992] = in_data[58015:57984] - in_data[58047:58016];
  assign out_data[29055:29024] = in_data[58079:58048] - in_data[58111:58080];
  assign out_data[29087:29056] = in_data[58143:58112] - in_data[58175:58144];
  assign out_data[2911:2880] = in_data[5791:5760] - in_data[5823:5792];
  assign out_data[29119:29088] = in_data[58207:58176] - in_data[58239:58208];
  assign out_data[29151:29120] = in_data[58271:58240] - in_data[58303:58272];
  assign out_data[29183:29152] = in_data[58335:58304] - in_data[58367:58336];
  assign out_data[29215:29184] = in_data[58399:58368] - in_data[58431:58400];
  assign out_data[29247:29216] = in_data[58463:58432] - in_data[58495:58464];
  assign out_data[29279:29248] = in_data[58527:58496] - in_data[58559:58528];
  assign out_data[29311:29280] = in_data[58591:58560] - in_data[58623:58592];
  assign out_data[29343:29312] = in_data[58655:58624] - in_data[58687:58656];
  assign out_data[29375:29344] = in_data[58719:58688] - in_data[58751:58720];
  assign out_data[29407:29376] = in_data[58783:58752] - in_data[58815:58784];
  assign out_data[2943:2912] = in_data[5855:5824] - in_data[5887:5856];
  assign out_data[29439:29408] = in_data[58847:58816] - in_data[58879:58848];
  assign out_data[29471:29440] = in_data[58911:58880] - in_data[58943:58912];
  assign out_data[29503:29472] = in_data[58975:58944] - in_data[59007:58976];
  assign out_data[29535:29504] = in_data[59039:59008] - in_data[59071:59040];
  assign out_data[29567:29536] = in_data[59103:59072] - in_data[59135:59104];
  assign out_data[29599:29568] = in_data[59167:59136] - in_data[59199:59168];
  assign out_data[29631:29600] = in_data[59231:59200] - in_data[59263:59232];
  assign out_data[29663:29632] = in_data[59295:59264] - in_data[59327:59296];
  assign out_data[29695:29664] = in_data[59359:59328] - in_data[59391:59360];
  assign out_data[29727:29696] = in_data[59423:59392] - in_data[59455:59424];
  assign out_data[2975:2944] = in_data[5919:5888] - in_data[5951:5920];
  assign out_data[29759:29728] = in_data[59487:59456] - in_data[59519:59488];
  assign out_data[29791:29760] = in_data[59551:59520] - in_data[59583:59552];
  assign out_data[29823:29792] = in_data[59615:59584] - in_data[59647:59616];
  assign out_data[29855:29824] = in_data[59679:59648] - in_data[59711:59680];
  assign out_data[29887:29856] = in_data[59743:59712] - in_data[59775:59744];
  assign out_data[29919:29888] = in_data[59807:59776] - in_data[59839:59808];
  assign out_data[29951:29920] = in_data[59871:59840] - in_data[59903:59872];
  assign out_data[29983:29952] = in_data[59935:59904] - in_data[59967:59936];
  assign out_data[30015:29984] = in_data[59999:59968] - in_data[60031:60000];
  assign out_data[30047:30016] = in_data[60063:60032] - in_data[60095:60064];
  assign out_data[3007:2976] = in_data[5983:5952] - in_data[6015:5984];
  assign out_data[30079:30048] = in_data[60127:60096] - in_data[60159:60128];
  assign out_data[30111:30080] = in_data[60191:60160] - in_data[60223:60192];
  assign out_data[30143:30112] = in_data[60255:60224] - in_data[60287:60256];
  assign out_data[30175:30144] = in_data[60319:60288] - in_data[60351:60320];
  assign out_data[30207:30176] = in_data[60383:60352] - in_data[60415:60384];
  assign out_data[30239:30208] = in_data[60447:60416] - in_data[60479:60448];
  assign out_data[30271:30240] = in_data[60511:60480] - in_data[60543:60512];
  assign out_data[30303:30272] = in_data[60575:60544] - in_data[60607:60576];
  assign out_data[30335:30304] = in_data[60639:60608] - in_data[60671:60640];
  assign out_data[30367:30336] = in_data[60703:60672] - in_data[60735:60704];
  assign out_data[3039:3008] = in_data[6047:6016] - in_data[6079:6048];
  assign out_data[30399:30368] = in_data[60767:60736] - in_data[60799:60768];
  assign out_data[30431:30400] = in_data[60831:60800] - in_data[60863:60832];
  assign out_data[30463:30432] = in_data[60895:60864] - in_data[60927:60896];
  assign out_data[30495:30464] = in_data[60959:60928] - in_data[60991:60960];
  assign out_data[30527:30496] = in_data[61023:60992] - in_data[61055:61024];
  assign out_data[30559:30528] = in_data[61087:61056] - in_data[61119:61088];
  assign out_data[30591:30560] = in_data[61151:61120] - in_data[61183:61152];
  assign out_data[30623:30592] = in_data[61215:61184] - in_data[61247:61216];
  assign out_data[30655:30624] = in_data[61279:61248] - in_data[61311:61280];
  assign out_data[30687:30656] = in_data[61343:61312] - in_data[61375:61344];
  assign out_data[3071:3040] = in_data[6111:6080] - in_data[6143:6112];
  assign out_data[30719:30688] = in_data[61407:61376] - in_data[61439:61408];
  assign out_data[30751:30720] = in_data[61471:61440] - in_data[61503:61472];
  assign out_data[30783:30752] = in_data[61535:61504] - in_data[61567:61536];
  assign out_data[30815:30784] = in_data[61599:61568] - in_data[61631:61600];
  assign out_data[30847:30816] = in_data[61663:61632] - in_data[61695:61664];
  assign out_data[30879:30848] = in_data[61727:61696] - in_data[61759:61728];
  assign out_data[30911:30880] = in_data[61791:61760] - in_data[61823:61792];
  assign out_data[30943:30912] = in_data[61855:61824] - in_data[61887:61856];
  assign out_data[30975:30944] = in_data[61919:61888] - in_data[61951:61920];
  assign out_data[31007:30976] = in_data[61983:61952] - in_data[62015:61984];
  assign out_data[3103:3072] = in_data[6175:6144] - in_data[6207:6176];
  assign out_data[31039:31008] = in_data[62047:62016] - in_data[62079:62048];
  assign out_data[31071:31040] = in_data[62111:62080] - in_data[62143:62112];
  assign out_data[31103:31072] = in_data[62175:62144] - in_data[62207:62176];
  assign out_data[31135:31104] = in_data[62239:62208] - in_data[62271:62240];
  assign out_data[31167:31136] = in_data[62303:62272] - in_data[62335:62304];
  assign out_data[31199:31168] = in_data[62367:62336] - in_data[62399:62368];
  assign out_data[31231:31200] = in_data[62431:62400] - in_data[62463:62432];
  assign out_data[31263:31232] = in_data[62495:62464] - in_data[62527:62496];
  assign out_data[31295:31264] = in_data[62559:62528] - in_data[62591:62560];
  assign out_data[31327:31296] = in_data[62623:62592] - in_data[62655:62624];
  assign out_data[3135:3104] = in_data[6239:6208] - in_data[6271:6240];
  assign out_data[31359:31328] = in_data[62687:62656] - in_data[62719:62688];
  assign out_data[31391:31360] = in_data[62751:62720] - in_data[62783:62752];
  assign out_data[31423:31392] = in_data[62815:62784] - in_data[62847:62816];
  assign out_data[31455:31424] = in_data[62879:62848] - in_data[62911:62880];
  assign out_data[31487:31456] = in_data[62943:62912] - in_data[62975:62944];
  assign out_data[31519:31488] = in_data[63007:62976] - in_data[63039:63008];
  assign out_data[31551:31520] = in_data[63071:63040] - in_data[63103:63072];
  assign out_data[31583:31552] = in_data[63135:63104] - in_data[63167:63136];
  assign out_data[31615:31584] = in_data[63199:63168] - in_data[63231:63200];
  assign out_data[31647:31616] = in_data[63263:63232] - in_data[63295:63264];
  assign out_data[3167:3136] = in_data[6303:6272] - in_data[6335:6304];
  assign out_data[31679:31648] = in_data[63327:63296] - in_data[63359:63328];
  assign out_data[31711:31680] = in_data[63391:63360] - in_data[63423:63392];
  assign out_data[31743:31712] = in_data[63455:63424] - in_data[63487:63456];
  assign out_data[31775:31744] = in_data[63519:63488] - in_data[63551:63520];
  assign out_data[31807:31776] = in_data[63583:63552] - in_data[63615:63584];
  assign out_data[31839:31808] = in_data[63647:63616] - in_data[63679:63648];
  assign out_data[31871:31840] = in_data[63711:63680] - in_data[63743:63712];
  assign out_data[31903:31872] = in_data[63775:63744] - in_data[63807:63776];
  assign out_data[31935:31904] = in_data[63839:63808] - in_data[63871:63840];
  assign out_data[31967:31936] = in_data[63903:63872] - in_data[63935:63904];
  assign out_data[31:0] = in_data[31:0] - in_data[63:32];
  assign out_data[319:288] = in_data[607:576] - in_data[639:608];
  assign out_data[3199:3168] = in_data[6367:6336] - in_data[6399:6368];
  assign out_data[31999:31968] = in_data[63967:63936] - in_data[63999:63968];
  assign out_data[32031:32000] = in_data[64031:64000] - in_data[64063:64032];
  assign out_data[32063:32032] = in_data[64095:64064] - in_data[64127:64096];
  assign out_data[32095:32064] = in_data[64159:64128] - in_data[64191:64160];
  assign out_data[32127:32096] = in_data[64223:64192] - in_data[64255:64224];
  assign out_data[32159:32128] = in_data[64287:64256] - in_data[64319:64288];
  assign out_data[32191:32160] = in_data[64351:64320] - in_data[64383:64352];
  assign out_data[32223:32192] = in_data[64415:64384] - in_data[64447:64416];
  assign out_data[32255:32224] = in_data[64479:64448] - in_data[64511:64480];
  assign out_data[32287:32256] = in_data[64543:64512] - in_data[64575:64544];
  assign out_data[3231:3200] = in_data[6431:6400] - in_data[6463:6432];
  assign out_data[32319:32288] = in_data[64607:64576] - in_data[64639:64608];
  assign out_data[32351:32320] = in_data[64671:64640] - in_data[64703:64672];
  assign out_data[32383:32352] = in_data[64735:64704] - in_data[64767:64736];
  assign out_data[32415:32384] = in_data[64799:64768] - in_data[64831:64800];
  assign out_data[32447:32416] = in_data[64863:64832] - in_data[64895:64864];
  assign out_data[32479:32448] = in_data[64927:64896] - in_data[64959:64928];
  assign out_data[32511:32480] = in_data[64991:64960] - in_data[65023:64992];
  assign out_data[32543:32512] = in_data[65055:65024] - in_data[65087:65056];
  assign out_data[32575:32544] = in_data[65119:65088] - in_data[65151:65120];
  assign out_data[32607:32576] = in_data[65183:65152] - in_data[65215:65184];
  assign out_data[3263:3232] = in_data[6495:6464] - in_data[6527:6496];
  assign out_data[32639:32608] = in_data[65247:65216] - in_data[65279:65248];
  assign out_data[32671:32640] = in_data[65311:65280] - in_data[65343:65312];
  assign out_data[32703:32672] = in_data[65375:65344] - in_data[65407:65376];
  assign out_data[32735:32704] = in_data[65439:65408] - in_data[65471:65440];
  assign out_data[32767:32736] = in_data[65503:65472] - in_data[65535:65504];
  assign out_data[32799:32768] = in_data[65567:65536] - in_data[65599:65568];
  assign out_data[32831:32800] = in_data[65631:65600] - in_data[65663:65632];
  assign out_data[32863:32832] = in_data[65695:65664] - in_data[65727:65696];
  assign out_data[32895:32864] = in_data[65759:65728] - in_data[65791:65760];
  assign out_data[32927:32896] = in_data[65823:65792] - in_data[65855:65824];
  assign out_data[3295:3264] = in_data[6559:6528] - in_data[6591:6560];
  assign out_data[32959:32928] = in_data[65887:65856] - in_data[65919:65888];
  assign out_data[32991:32960] = in_data[65951:65920] - in_data[65983:65952];
  assign out_data[33023:32992] = in_data[66015:65984] - in_data[66047:66016];
  assign out_data[33055:33024] = in_data[66079:66048] - in_data[66111:66080];
  assign out_data[33087:33056] = in_data[66143:66112] - in_data[66175:66144];
  assign out_data[33119:33088] = in_data[66207:66176] - in_data[66239:66208];
  assign out_data[33151:33120] = in_data[66271:66240] - in_data[66303:66272];
  assign out_data[33183:33152] = in_data[66335:66304] - in_data[66367:66336];
  assign out_data[33215:33184] = in_data[66399:66368] - in_data[66431:66400];
  assign out_data[33247:33216] = in_data[66463:66432] - in_data[66495:66464];
  assign out_data[3327:3296] = in_data[6623:6592] - in_data[6655:6624];
  assign out_data[33279:33248] = in_data[66527:66496] - in_data[66559:66528];
  assign out_data[33311:33280] = in_data[66591:66560] - in_data[66623:66592];
  assign out_data[33343:33312] = in_data[66655:66624] - in_data[66687:66656];
  assign out_data[33375:33344] = in_data[66719:66688] - in_data[66751:66720];
  assign out_data[33407:33376] = in_data[66783:66752] - in_data[66815:66784];
  assign out_data[33439:33408] = in_data[66847:66816] - in_data[66879:66848];
  assign out_data[33471:33440] = in_data[66911:66880] - in_data[66943:66912];
  assign out_data[33503:33472] = in_data[66975:66944] - in_data[67007:66976];
  assign out_data[33535:33504] = in_data[67039:67008] - in_data[67071:67040];
  assign out_data[33567:33536] = in_data[67103:67072] - in_data[67135:67104];
  assign out_data[3359:3328] = in_data[6687:6656] - in_data[6719:6688];
  assign out_data[33599:33568] = in_data[67167:67136] - in_data[67199:67168];
  assign out_data[33631:33600] = in_data[67231:67200] - in_data[67263:67232];
  assign out_data[33663:33632] = in_data[67295:67264] - in_data[67327:67296];
  assign out_data[33695:33664] = in_data[67359:67328] - in_data[67391:67360];
  assign out_data[33727:33696] = in_data[67423:67392] - in_data[67455:67424];
  assign out_data[33759:33728] = in_data[67487:67456] - in_data[67519:67488];
  assign out_data[33791:33760] = in_data[67551:67520] - in_data[67583:67552];
  assign out_data[33823:33792] = in_data[67615:67584] - in_data[67647:67616];
  assign out_data[33855:33824] = in_data[67679:67648] - in_data[67711:67680];
  assign out_data[33887:33856] = in_data[67743:67712] - in_data[67775:67744];
  assign out_data[3391:3360] = in_data[6751:6720] - in_data[6783:6752];
  assign out_data[33919:33888] = in_data[67807:67776] - in_data[67839:67808];
  assign out_data[33951:33920] = in_data[67871:67840] - in_data[67903:67872];
  assign out_data[33983:33952] = in_data[67935:67904] - in_data[67967:67936];
  assign out_data[34015:33984] = in_data[67999:67968] - in_data[68031:68000];
  assign out_data[34047:34016] = in_data[68063:68032] - in_data[68095:68064];
  assign out_data[34079:34048] = in_data[68127:68096] - in_data[68159:68128];
  assign out_data[34111:34080] = in_data[68191:68160] - in_data[68223:68192];
  assign out_data[34143:34112] = in_data[68255:68224] - in_data[68287:68256];
  assign out_data[34175:34144] = in_data[68319:68288] - in_data[68351:68320];
  assign out_data[34207:34176] = in_data[68383:68352] - in_data[68415:68384];
  assign out_data[3423:3392] = in_data[6815:6784] - in_data[6847:6816];
  assign out_data[34239:34208] = in_data[68447:68416] - in_data[68479:68448];
  assign out_data[34271:34240] = in_data[68511:68480] - in_data[68543:68512];
  assign out_data[34303:34272] = in_data[68575:68544] - in_data[68607:68576];
  assign out_data[34335:34304] = in_data[68639:68608] - in_data[68671:68640];
  assign out_data[34367:34336] = in_data[68703:68672] - in_data[68735:68704];
  assign out_data[34399:34368] = in_data[68767:68736] - in_data[68799:68768];
  assign out_data[34431:34400] = in_data[68831:68800] - in_data[68863:68832];
  assign out_data[34463:34432] = in_data[68895:68864] - in_data[68927:68896];
  assign out_data[34495:34464] = in_data[68959:68928] - in_data[68991:68960];
  assign out_data[34527:34496] = in_data[69023:68992] - in_data[69055:69024];
  assign out_data[3455:3424] = in_data[6879:6848] - in_data[6911:6880];
  assign out_data[34559:34528] = in_data[69087:69056] - in_data[69119:69088];
  assign out_data[34591:34560] = in_data[69151:69120] - in_data[69183:69152];
  assign out_data[34623:34592] = in_data[69215:69184] - in_data[69247:69216];
  assign out_data[34655:34624] = in_data[69279:69248] - in_data[69311:69280];
  assign out_data[34687:34656] = in_data[69343:69312] - in_data[69375:69344];
  assign out_data[34719:34688] = in_data[69407:69376] - in_data[69439:69408];
  assign out_data[34751:34720] = in_data[69471:69440] - in_data[69503:69472];
  assign out_data[34783:34752] = in_data[69535:69504] - in_data[69567:69536];
  assign out_data[34815:34784] = in_data[69599:69568] - in_data[69631:69600];
  assign out_data[34847:34816] = in_data[69663:69632] - in_data[69695:69664];
  assign out_data[3487:3456] = in_data[6943:6912] - in_data[6975:6944];
  assign out_data[34879:34848] = in_data[69727:69696] - in_data[69759:69728];
  assign out_data[34911:34880] = in_data[69791:69760] - in_data[69823:69792];
  assign out_data[34943:34912] = in_data[69855:69824] - in_data[69887:69856];
  assign out_data[34975:34944] = in_data[69919:69888] - in_data[69951:69920];
  assign out_data[35007:34976] = in_data[69983:69952] - in_data[70015:69984];
  assign out_data[35039:35008] = in_data[70047:70016] - in_data[70079:70048];
  assign out_data[35071:35040] = in_data[70111:70080] - in_data[70143:70112];
  assign out_data[35103:35072] = in_data[70175:70144] - in_data[70207:70176];
  assign out_data[35135:35104] = in_data[70239:70208] - in_data[70271:70240];
  assign out_data[35167:35136] = in_data[70303:70272] - in_data[70335:70304];
  assign out_data[351:320] = in_data[671:640] - in_data[703:672];
  assign out_data[3519:3488] = in_data[7007:6976] - in_data[7039:7008];
  assign out_data[35199:35168] = in_data[70367:70336] - in_data[70399:70368];
  assign out_data[35231:35200] = in_data[70431:70400] - in_data[70463:70432];
  assign out_data[35263:35232] = in_data[70495:70464] - in_data[70527:70496];
  assign out_data[35295:35264] = in_data[70559:70528] - in_data[70591:70560];
  assign out_data[35327:35296] = in_data[70623:70592] - in_data[70655:70624];
  assign out_data[35359:35328] = in_data[70687:70656] - in_data[70719:70688];
  assign out_data[35391:35360] = in_data[70751:70720] - in_data[70783:70752];
  assign out_data[35423:35392] = in_data[70815:70784] - in_data[70847:70816];
  assign out_data[35455:35424] = in_data[70879:70848] - in_data[70911:70880];
  assign out_data[35487:35456] = in_data[70943:70912] - in_data[70975:70944];
  assign out_data[3551:3520] = in_data[7071:7040] - in_data[7103:7072];
  assign out_data[35519:35488] = in_data[71007:70976] - in_data[71039:71008];
  assign out_data[35551:35520] = in_data[71071:71040] - in_data[71103:71072];
  assign out_data[35583:35552] = in_data[71135:71104] - in_data[71167:71136];
  assign out_data[35615:35584] = in_data[71199:71168] - in_data[71231:71200];
  assign out_data[35647:35616] = in_data[71263:71232] - in_data[71295:71264];
  assign out_data[35679:35648] = in_data[71327:71296] - in_data[71359:71328];
  assign out_data[35711:35680] = in_data[71391:71360] - in_data[71423:71392];
  assign out_data[35743:35712] = in_data[71455:71424] - in_data[71487:71456];
  assign out_data[35775:35744] = in_data[71519:71488] - in_data[71551:71520];
  assign out_data[35807:35776] = in_data[71583:71552] - in_data[71615:71584];
  assign out_data[3583:3552] = in_data[7135:7104] - in_data[7167:7136];
  assign out_data[35839:35808] = in_data[71647:71616] - in_data[71679:71648];
  assign out_data[35871:35840] = in_data[71711:71680] - in_data[71743:71712];
  assign out_data[35903:35872] = in_data[71775:71744] - in_data[71807:71776];
  assign out_data[35935:35904] = in_data[71839:71808] - in_data[71871:71840];
  assign out_data[35967:35936] = in_data[71903:71872] - in_data[71935:71904];
  assign out_data[35999:35968] = in_data[71967:71936] - in_data[71999:71968];
  assign out_data[36031:36000] = in_data[72031:72000] - in_data[72063:72032];
  assign out_data[36063:36032] = in_data[72095:72064] - in_data[72127:72096];
  assign out_data[36095:36064] = in_data[72159:72128] - in_data[72191:72160];
  assign out_data[36127:36096] = in_data[72223:72192] - in_data[72255:72224];
  assign out_data[3615:3584] = in_data[7199:7168] - in_data[7231:7200];
  assign out_data[36159:36128] = in_data[72287:72256] - in_data[72319:72288];
  assign out_data[36191:36160] = in_data[72351:72320] - in_data[72383:72352];
  assign out_data[36223:36192] = in_data[72415:72384] - in_data[72447:72416];
  assign out_data[36255:36224] = in_data[72479:72448] - in_data[72511:72480];
  assign out_data[36287:36256] = in_data[72543:72512] - in_data[72575:72544];
  assign out_data[36319:36288] = in_data[72607:72576] - in_data[72639:72608];
  assign out_data[36351:36320] = in_data[72671:72640] - in_data[72703:72672];
  assign out_data[36383:36352] = in_data[72735:72704] - in_data[72767:72736];
  assign out_data[36415:36384] = in_data[72799:72768] - in_data[72831:72800];
  assign out_data[36447:36416] = in_data[72863:72832] - in_data[72895:72864];
  assign out_data[3647:3616] = in_data[7263:7232] - in_data[7295:7264];
  assign out_data[36479:36448] = in_data[72927:72896] - in_data[72959:72928];
  assign out_data[36511:36480] = in_data[72991:72960] - in_data[73023:72992];
  assign out_data[36543:36512] = in_data[73055:73024] - in_data[73087:73056];
  assign out_data[36575:36544] = in_data[73119:73088] - in_data[73151:73120];
  assign out_data[36607:36576] = in_data[73183:73152] - in_data[73215:73184];
  assign out_data[36639:36608] = in_data[73247:73216] - in_data[73279:73248];
  assign out_data[36671:36640] = in_data[73311:73280] - in_data[73343:73312];
  assign out_data[36703:36672] = in_data[73375:73344] - in_data[73407:73376];
  assign out_data[36735:36704] = in_data[73439:73408] - in_data[73471:73440];
  assign out_data[36767:36736] = in_data[73503:73472] - in_data[73535:73504];
  assign out_data[3679:3648] = in_data[7327:7296] - in_data[7359:7328];
  assign out_data[36799:36768] = in_data[73567:73536] - in_data[73599:73568];
  assign out_data[36831:36800] = in_data[73631:73600] - in_data[73663:73632];
  assign out_data[36863:36832] = in_data[73695:73664] - in_data[73727:73696];
  assign out_data[36895:36864] = in_data[73759:73728] - in_data[73791:73760];
  assign out_data[36927:36896] = in_data[73823:73792] - in_data[73855:73824];
  assign out_data[36959:36928] = in_data[73887:73856] - in_data[73919:73888];
  assign out_data[36991:36960] = in_data[73951:73920] - in_data[73983:73952];
  assign out_data[37023:36992] = in_data[74015:73984] - in_data[74047:74016];
  assign out_data[37055:37024] = in_data[74079:74048] - in_data[74111:74080];
  assign out_data[37087:37056] = in_data[74143:74112] - in_data[74175:74144];
  assign out_data[3711:3680] = in_data[7391:7360] - in_data[7423:7392];
  assign out_data[37119:37088] = in_data[74207:74176] - in_data[74239:74208];
  assign out_data[37151:37120] = in_data[74271:74240] - in_data[74303:74272];
  assign out_data[37183:37152] = in_data[74335:74304] - in_data[74367:74336];
  assign out_data[37215:37184] = in_data[74399:74368] - in_data[74431:74400];
  assign out_data[37247:37216] = in_data[74463:74432] - in_data[74495:74464];
  assign out_data[37279:37248] = in_data[74527:74496] - in_data[74559:74528];
  assign out_data[37311:37280] = in_data[74591:74560] - in_data[74623:74592];
  assign out_data[37343:37312] = in_data[74655:74624] - in_data[74687:74656];
  assign out_data[37375:37344] = in_data[74719:74688] - in_data[74751:74720];
  assign out_data[37407:37376] = in_data[74783:74752] - in_data[74815:74784];
  assign out_data[3743:3712] = in_data[7455:7424] - in_data[7487:7456];
  assign out_data[37439:37408] = in_data[74847:74816] - in_data[74879:74848];
  assign out_data[37471:37440] = in_data[74911:74880] - in_data[74943:74912];
  assign out_data[37503:37472] = in_data[74975:74944] - in_data[75007:74976];
  assign out_data[37535:37504] = in_data[75039:75008] - in_data[75071:75040];
  assign out_data[37567:37536] = in_data[75103:75072] - in_data[75135:75104];
  assign out_data[37599:37568] = in_data[75167:75136] - in_data[75199:75168];
  assign out_data[37631:37600] = in_data[75231:75200] - in_data[75263:75232];
  assign out_data[37663:37632] = in_data[75295:75264] - in_data[75327:75296];
  assign out_data[37695:37664] = in_data[75359:75328] - in_data[75391:75360];
  assign out_data[37727:37696] = in_data[75423:75392] - in_data[75455:75424];
  assign out_data[3775:3744] = in_data[7519:7488] - in_data[7551:7520];
  assign out_data[37759:37728] = in_data[75487:75456] - in_data[75519:75488];
  assign out_data[37791:37760] = in_data[75551:75520] - in_data[75583:75552];
  assign out_data[37823:37792] = in_data[75615:75584] - in_data[75647:75616];
  assign out_data[37855:37824] = in_data[75679:75648] - in_data[75711:75680];
  assign out_data[37887:37856] = in_data[75743:75712] - in_data[75775:75744];
  assign out_data[37919:37888] = in_data[75807:75776] - in_data[75839:75808];
  assign out_data[37951:37920] = in_data[75871:75840] - in_data[75903:75872];
  assign out_data[37983:37952] = in_data[75935:75904] - in_data[75967:75936];
  assign out_data[38015:37984] = in_data[75999:75968] - in_data[76031:76000];
  assign out_data[38047:38016] = in_data[76063:76032] - in_data[76095:76064];
  assign out_data[3807:3776] = in_data[7583:7552] - in_data[7615:7584];
  assign out_data[38079:38048] = in_data[76127:76096] - in_data[76159:76128];
  assign out_data[38111:38080] = in_data[76191:76160] - in_data[76223:76192];
  assign out_data[38143:38112] = in_data[76255:76224] - in_data[76287:76256];
  assign out_data[38175:38144] = in_data[76319:76288] - in_data[76351:76320];
  assign out_data[38207:38176] = in_data[76383:76352] - in_data[76415:76384];
  assign out_data[38239:38208] = in_data[76447:76416] - in_data[76479:76448];
  assign out_data[38271:38240] = in_data[76511:76480] - in_data[76543:76512];
  assign out_data[38303:38272] = in_data[76575:76544] - in_data[76607:76576];
  assign out_data[38335:38304] = in_data[76639:76608] - in_data[76671:76640];
  assign out_data[38367:38336] = in_data[76703:76672] - in_data[76735:76704];
  assign out_data[383:352] = in_data[735:704] - in_data[767:736];
  assign out_data[3839:3808] = in_data[7647:7616] - in_data[7679:7648];
  assign out_data[38399:38368] = in_data[76767:76736] - in_data[76799:76768];
  assign out_data[38431:38400] = in_data[76831:76800] - in_data[76863:76832];
  assign out_data[38463:38432] = in_data[76895:76864] - in_data[76927:76896];
  assign out_data[38495:38464] = in_data[76959:76928] - in_data[76991:76960];
  assign out_data[38527:38496] = in_data[77023:76992] - in_data[77055:77024];
  assign out_data[38559:38528] = in_data[77087:77056] - in_data[77119:77088];
  assign out_data[38591:38560] = in_data[77151:77120] - in_data[77183:77152];
  assign out_data[38623:38592] = in_data[77215:77184] - in_data[77247:77216];
  assign out_data[38655:38624] = in_data[77279:77248] - in_data[77311:77280];
  assign out_data[38687:38656] = in_data[77343:77312] - in_data[77375:77344];
  assign out_data[3871:3840] = in_data[7711:7680] - in_data[7743:7712];
  assign out_data[38719:38688] = in_data[77407:77376] - in_data[77439:77408];
  assign out_data[38751:38720] = in_data[77471:77440] - in_data[77503:77472];
  assign out_data[38783:38752] = in_data[77535:77504] - in_data[77567:77536];
  assign out_data[38815:38784] = in_data[77599:77568] - in_data[77631:77600];
  assign out_data[38847:38816] = in_data[77663:77632] - in_data[77695:77664];
  assign out_data[38879:38848] = in_data[77727:77696] - in_data[77759:77728];
  assign out_data[38911:38880] = in_data[77791:77760] - in_data[77823:77792];
  assign out_data[38943:38912] = in_data[77855:77824] - in_data[77887:77856];
  assign out_data[38975:38944] = in_data[77919:77888] - in_data[77951:77920];
  assign out_data[39007:38976] = in_data[77983:77952] - in_data[78015:77984];
  assign out_data[3903:3872] = in_data[7775:7744] - in_data[7807:7776];
  assign out_data[39039:39008] = in_data[78047:78016] - in_data[78079:78048];
  assign out_data[39071:39040] = in_data[78111:78080] - in_data[78143:78112];
  assign out_data[39103:39072] = in_data[78175:78144] - in_data[78207:78176];
  assign out_data[39135:39104] = in_data[78239:78208] - in_data[78271:78240];
  assign out_data[39167:39136] = in_data[78303:78272] - in_data[78335:78304];
  assign out_data[39199:39168] = in_data[78367:78336] - in_data[78399:78368];
  assign out_data[39231:39200] = in_data[78431:78400] - in_data[78463:78432];
  assign out_data[39263:39232] = in_data[78495:78464] - in_data[78527:78496];
  assign out_data[39295:39264] = in_data[78559:78528] - in_data[78591:78560];
  assign out_data[39327:39296] = in_data[78623:78592] - in_data[78655:78624];
  assign out_data[3935:3904] = in_data[7839:7808] - in_data[7871:7840];
  assign out_data[39359:39328] = in_data[78687:78656] - in_data[78719:78688];
  assign out_data[39391:39360] = in_data[78751:78720] - in_data[78783:78752];
  assign out_data[39423:39392] = in_data[78815:78784] - in_data[78847:78816];
  assign out_data[39455:39424] = in_data[78879:78848] - in_data[78911:78880];
  assign out_data[39487:39456] = in_data[78943:78912] - in_data[78975:78944];
  assign out_data[39519:39488] = in_data[79007:78976] - in_data[79039:79008];
  assign out_data[39551:39520] = in_data[79071:79040] - in_data[79103:79072];
  assign out_data[39583:39552] = in_data[79135:79104] - in_data[79167:79136];
  assign out_data[39615:39584] = in_data[79199:79168] - in_data[79231:79200];
  assign out_data[39647:39616] = in_data[79263:79232] - in_data[79295:79264];
  assign out_data[3967:3936] = in_data[7903:7872] - in_data[7935:7904];
  assign out_data[39679:39648] = in_data[79327:79296] - in_data[79359:79328];
  assign out_data[39711:39680] = in_data[79391:79360] - in_data[79423:79392];
  assign out_data[39743:39712] = in_data[79455:79424] - in_data[79487:79456];
  assign out_data[39775:39744] = in_data[79519:79488] - in_data[79551:79520];
  assign out_data[39807:39776] = in_data[79583:79552] - in_data[79615:79584];
  assign out_data[39839:39808] = in_data[79647:79616] - in_data[79679:79648];
  assign out_data[39871:39840] = in_data[79711:79680] - in_data[79743:79712];
  assign out_data[39903:39872] = in_data[79775:79744] - in_data[79807:79776];
  assign out_data[39935:39904] = in_data[79839:79808] - in_data[79871:79840];
  assign out_data[39967:39936] = in_data[79903:79872] - in_data[79935:79904];
  assign out_data[3999:3968] = in_data[7967:7936] - in_data[7999:7968];
  assign out_data[39999:39968] = in_data[79967:79936] - in_data[79999:79968];
  assign out_data[40031:40000] = in_data[80031:80000] - in_data[80063:80032];
  assign out_data[40063:40032] = in_data[80095:80064] - in_data[80127:80096];
  assign out_data[40095:40064] = in_data[80159:80128] - in_data[80191:80160];
  assign out_data[40127:40096] = in_data[80223:80192] - in_data[80255:80224];
  assign out_data[40159:40128] = in_data[80287:80256] - in_data[80319:80288];
  assign out_data[40191:40160] = in_data[80351:80320] - in_data[80383:80352];
  assign out_data[40223:40192] = in_data[80415:80384] - in_data[80447:80416];
  assign out_data[40255:40224] = in_data[80479:80448] - in_data[80511:80480];
  assign out_data[40287:40256] = in_data[80543:80512] - in_data[80575:80544];
  assign out_data[4031:4000] = in_data[8031:8000] - in_data[8063:8032];
  assign out_data[40319:40288] = in_data[80607:80576] - in_data[80639:80608];
  assign out_data[40351:40320] = in_data[80671:80640] - in_data[80703:80672];
  assign out_data[40383:40352] = in_data[80735:80704] - in_data[80767:80736];
  assign out_data[40415:40384] = in_data[80799:80768] - in_data[80831:80800];
  assign out_data[40447:40416] = in_data[80863:80832] - in_data[80895:80864];
  assign out_data[40479:40448] = in_data[80927:80896] - in_data[80959:80928];
  assign out_data[40511:40480] = in_data[80991:80960] - in_data[81023:80992];
  assign out_data[40543:40512] = in_data[81055:81024] - in_data[81087:81056];
  assign out_data[40575:40544] = in_data[81119:81088] - in_data[81151:81120];
  assign out_data[40607:40576] = in_data[81183:81152] - in_data[81215:81184];
  assign out_data[4063:4032] = in_data[8095:8064] - in_data[8127:8096];
  assign out_data[40639:40608] = in_data[81247:81216] - in_data[81279:81248];
  assign out_data[40671:40640] = in_data[81311:81280] - in_data[81343:81312];
  assign out_data[40703:40672] = in_data[81375:81344] - in_data[81407:81376];
  assign out_data[40735:40704] = in_data[81439:81408] - in_data[81471:81440];
  assign out_data[40767:40736] = in_data[81503:81472] - in_data[81535:81504];
  assign out_data[40799:40768] = in_data[81567:81536] - in_data[81599:81568];
  assign out_data[40831:40800] = in_data[81631:81600] - in_data[81663:81632];
  assign out_data[40863:40832] = in_data[81695:81664] - in_data[81727:81696];
  assign out_data[40895:40864] = in_data[81759:81728] - in_data[81791:81760];
  assign out_data[40927:40896] = in_data[81823:81792] - in_data[81855:81824];
  assign out_data[4095:4064] = in_data[8159:8128] - in_data[8191:8160];
  assign out_data[40959:40928] = in_data[81887:81856] - in_data[81919:81888];
  assign out_data[40991:40960] = in_data[81951:81920] - in_data[81983:81952];
  assign out_data[41023:40992] = in_data[82015:81984] - in_data[82047:82016];
  assign out_data[41055:41024] = in_data[82079:82048] - in_data[82111:82080];
  assign out_data[41087:41056] = in_data[82143:82112] - in_data[82175:82144];
  assign out_data[41119:41088] = in_data[82207:82176] - in_data[82239:82208];
  assign out_data[41151:41120] = in_data[82271:82240] - in_data[82303:82272];
  assign out_data[41183:41152] = in_data[82335:82304] - in_data[82367:82336];
  assign out_data[41215:41184] = in_data[82399:82368] - in_data[82431:82400];
  assign out_data[41247:41216] = in_data[82463:82432] - in_data[82495:82464];
  assign out_data[4127:4096] = in_data[8223:8192] - in_data[8255:8224];
  assign out_data[41279:41248] = in_data[82527:82496] - in_data[82559:82528];
  assign out_data[41311:41280] = in_data[82591:82560] - in_data[82623:82592];
  assign out_data[41343:41312] = in_data[82655:82624] - in_data[82687:82656];
  assign out_data[41375:41344] = in_data[82719:82688] - in_data[82751:82720];
  assign out_data[41407:41376] = in_data[82783:82752] - in_data[82815:82784];
  assign out_data[41439:41408] = in_data[82847:82816] - in_data[82879:82848];
  assign out_data[41471:41440] = in_data[82911:82880] - in_data[82943:82912];
  assign out_data[41503:41472] = in_data[82975:82944] - in_data[83007:82976];
  assign out_data[41535:41504] = in_data[83039:83008] - in_data[83071:83040];
  assign out_data[41567:41536] = in_data[83103:83072] - in_data[83135:83104];
  assign out_data[415:384] = in_data[799:768] - in_data[831:800];
  assign out_data[4159:4128] = in_data[8287:8256] - in_data[8319:8288];
  assign out_data[41599:41568] = in_data[83167:83136] - in_data[83199:83168];
  assign out_data[41631:41600] = in_data[83231:83200] - in_data[83263:83232];
  assign out_data[41663:41632] = in_data[83295:83264] - in_data[83327:83296];
  assign out_data[41695:41664] = in_data[83359:83328] - in_data[83391:83360];
  assign out_data[41727:41696] = in_data[83423:83392] - in_data[83455:83424];
  assign out_data[41759:41728] = in_data[83487:83456] - in_data[83519:83488];
  assign out_data[41791:41760] = in_data[83551:83520] - in_data[83583:83552];
  assign out_data[41823:41792] = in_data[83615:83584] - in_data[83647:83616];
  assign out_data[41855:41824] = in_data[83679:83648] - in_data[83711:83680];
  assign out_data[41887:41856] = in_data[83743:83712] - in_data[83775:83744];
  assign out_data[4191:4160] = in_data[8351:8320] - in_data[8383:8352];
  assign out_data[41919:41888] = in_data[83807:83776] - in_data[83839:83808];
  assign out_data[41951:41920] = in_data[83871:83840] - in_data[83903:83872];
  assign out_data[41983:41952] = in_data[83935:83904] - in_data[83967:83936];
  assign out_data[42015:41984] = in_data[83999:83968] - in_data[84031:84000];
  assign out_data[42047:42016] = in_data[84063:84032] - in_data[84095:84064];
  assign out_data[42079:42048] = in_data[84127:84096] - in_data[84159:84128];
  assign out_data[42111:42080] = in_data[84191:84160] - in_data[84223:84192];
  assign out_data[42143:42112] = in_data[84255:84224] - in_data[84287:84256];
  assign out_data[42175:42144] = in_data[84319:84288] - in_data[84351:84320];
  assign out_data[42207:42176] = in_data[84383:84352] - in_data[84415:84384];
  assign out_data[4223:4192] = in_data[8415:8384] - in_data[8447:8416];
  assign out_data[42239:42208] = in_data[84447:84416] - in_data[84479:84448];
  assign out_data[42271:42240] = in_data[84511:84480] - in_data[84543:84512];
  assign out_data[42303:42272] = in_data[84575:84544] - in_data[84607:84576];
  assign out_data[42335:42304] = in_data[84639:84608] - in_data[84671:84640];
  assign out_data[42367:42336] = in_data[84703:84672] - in_data[84735:84704];
  assign out_data[42399:42368] = in_data[84767:84736] - in_data[84799:84768];
  assign out_data[42431:42400] = in_data[84831:84800] - in_data[84863:84832];
  assign out_data[42463:42432] = in_data[84895:84864] - in_data[84927:84896];
  assign out_data[42495:42464] = in_data[84959:84928] - in_data[84991:84960];
  assign out_data[42527:42496] = in_data[85023:84992] - in_data[85055:85024];
  assign out_data[4255:4224] = in_data[8479:8448] - in_data[8511:8480];
  assign out_data[42559:42528] = in_data[85087:85056] - in_data[85119:85088];
  assign out_data[42591:42560] = in_data[85151:85120] - in_data[85183:85152];
  assign out_data[42623:42592] = in_data[85215:85184] - in_data[85247:85216];
  assign out_data[42655:42624] = in_data[85279:85248] - in_data[85311:85280];
  assign out_data[42687:42656] = in_data[85343:85312] - in_data[85375:85344];
  assign out_data[42719:42688] = in_data[85407:85376] - in_data[85439:85408];
  assign out_data[42751:42720] = in_data[85471:85440] - in_data[85503:85472];
  assign out_data[42783:42752] = in_data[85535:85504] - in_data[85567:85536];
  assign out_data[42815:42784] = in_data[85599:85568] - in_data[85631:85600];
  assign out_data[42847:42816] = in_data[85663:85632] - in_data[85695:85664];
  assign out_data[4287:4256] = in_data[8543:8512] - in_data[8575:8544];
  assign out_data[42879:42848] = in_data[85727:85696] - in_data[85759:85728];
  assign out_data[42911:42880] = in_data[85791:85760] - in_data[85823:85792];
  assign out_data[42943:42912] = in_data[85855:85824] - in_data[85887:85856];
  assign out_data[42975:42944] = in_data[85919:85888] - in_data[85951:85920];
  assign out_data[43007:42976] = in_data[85983:85952] - in_data[86015:85984];
  assign out_data[43039:43008] = in_data[86047:86016] - in_data[86079:86048];
  assign out_data[43071:43040] = in_data[86111:86080] - in_data[86143:86112];
  assign out_data[43103:43072] = in_data[86175:86144] - in_data[86207:86176];
  assign out_data[43135:43104] = in_data[86239:86208] - in_data[86271:86240];
  assign out_data[43167:43136] = in_data[86303:86272] - in_data[86335:86304];
  assign out_data[4319:4288] = in_data[8607:8576] - in_data[8639:8608];
  assign out_data[43199:43168] = in_data[86367:86336] - in_data[86399:86368];
  assign out_data[43231:43200] = in_data[86431:86400] - in_data[86463:86432];
  assign out_data[43263:43232] = in_data[86495:86464] - in_data[86527:86496];
  assign out_data[43295:43264] = in_data[86559:86528] - in_data[86591:86560];
  assign out_data[43327:43296] = in_data[86623:86592] - in_data[86655:86624];
  assign out_data[43359:43328] = in_data[86687:86656] - in_data[86719:86688];
  assign out_data[43391:43360] = in_data[86751:86720] - in_data[86783:86752];
  assign out_data[43423:43392] = in_data[86815:86784] - in_data[86847:86816];
  assign out_data[43455:43424] = in_data[86879:86848] - in_data[86911:86880];
  assign out_data[43487:43456] = in_data[86943:86912] - in_data[86975:86944];
  assign out_data[4351:4320] = in_data[8671:8640] - in_data[8703:8672];
  assign out_data[43519:43488] = in_data[87007:86976] - in_data[87039:87008];
  assign out_data[43551:43520] = in_data[87071:87040] - in_data[87103:87072];
  assign out_data[43583:43552] = in_data[87135:87104] - in_data[87167:87136];
  assign out_data[43615:43584] = in_data[87199:87168] - in_data[87231:87200];
  assign out_data[43647:43616] = in_data[87263:87232] - in_data[87295:87264];
  assign out_data[43679:43648] = in_data[87327:87296] - in_data[87359:87328];
  assign out_data[43711:43680] = in_data[87391:87360] - in_data[87423:87392];
  assign out_data[43743:43712] = in_data[87455:87424] - in_data[87487:87456];
  assign out_data[43775:43744] = in_data[87519:87488] - in_data[87551:87520];
  assign out_data[43807:43776] = in_data[87583:87552] - in_data[87615:87584];
  assign out_data[4383:4352] = in_data[8735:8704] - in_data[8767:8736];
  assign out_data[43839:43808] = in_data[87647:87616] - in_data[87679:87648];
  assign out_data[43871:43840] = in_data[87711:87680] - in_data[87743:87712];
  assign out_data[43903:43872] = in_data[87775:87744] - in_data[87807:87776];
  assign out_data[43935:43904] = in_data[87839:87808] - in_data[87871:87840];
  assign out_data[43967:43936] = in_data[87903:87872] - in_data[87935:87904];
  assign out_data[43999:43968] = in_data[87967:87936] - in_data[87999:87968];
  assign out_data[44031:44000] = in_data[88031:88000] - in_data[88063:88032];
  assign out_data[44063:44032] = in_data[88095:88064] - in_data[88127:88096];
  assign out_data[44095:44064] = in_data[88159:88128] - in_data[88191:88160];
  assign out_data[44127:44096] = in_data[88223:88192] - in_data[88255:88224];
  assign out_data[4415:4384] = in_data[8799:8768] - in_data[8831:8800];
  assign out_data[44159:44128] = in_data[88287:88256] - in_data[88319:88288];
  assign out_data[44191:44160] = in_data[88351:88320] - in_data[88383:88352];
  assign out_data[44223:44192] = in_data[88415:88384] - in_data[88447:88416];
  assign out_data[44255:44224] = in_data[88479:88448] - in_data[88511:88480];
  assign out_data[44287:44256] = in_data[88543:88512] - in_data[88575:88544];
  assign out_data[44319:44288] = in_data[88607:88576] - in_data[88639:88608];
  assign out_data[44351:44320] = in_data[88671:88640] - in_data[88703:88672];
  assign out_data[44383:44352] = in_data[88735:88704] - in_data[88767:88736];
  assign out_data[44415:44384] = in_data[88799:88768] - in_data[88831:88800];
  assign out_data[44447:44416] = in_data[88863:88832] - in_data[88895:88864];
  assign out_data[4447:4416] = in_data[8863:8832] - in_data[8895:8864];
  assign out_data[44479:44448] = in_data[88927:88896] - in_data[88959:88928];
  assign out_data[44511:44480] = in_data[88991:88960] - in_data[89023:88992];
  assign out_data[44543:44512] = in_data[89055:89024] - in_data[89087:89056];
  assign out_data[44575:44544] = in_data[89119:89088] - in_data[89151:89120];
  assign out_data[44607:44576] = in_data[89183:89152] - in_data[89215:89184];
  assign out_data[44639:44608] = in_data[89247:89216] - in_data[89279:89248];
  assign out_data[44671:44640] = in_data[89311:89280] - in_data[89343:89312];
  assign out_data[44703:44672] = in_data[89375:89344] - in_data[89407:89376];
  assign out_data[44735:44704] = in_data[89439:89408] - in_data[89471:89440];
  assign out_data[44767:44736] = in_data[89503:89472] - in_data[89535:89504];
  assign out_data[447:416] = in_data[863:832] - in_data[895:864];
  assign out_data[4479:4448] = in_data[8927:8896] - in_data[8959:8928];
  assign out_data[44799:44768] = in_data[89567:89536] - in_data[89599:89568];
  assign out_data[44831:44800] = in_data[89631:89600] - in_data[89663:89632];
  assign out_data[44863:44832] = in_data[89695:89664] - in_data[89727:89696];
  assign out_data[44895:44864] = in_data[89759:89728] - in_data[89791:89760];
  assign out_data[44927:44896] = in_data[89823:89792] - in_data[89855:89824];
  assign out_data[44959:44928] = in_data[89887:89856] - in_data[89919:89888];
  assign out_data[44991:44960] = in_data[89951:89920] - in_data[89983:89952];
  assign out_data[45023:44992] = in_data[90015:89984] - in_data[90047:90016];
  assign out_data[45055:45024] = in_data[90079:90048] - in_data[90111:90080];
  assign out_data[45087:45056] = in_data[90143:90112] - in_data[90175:90144];
  assign out_data[4511:4480] = in_data[8991:8960] - in_data[9023:8992];
  assign out_data[45119:45088] = in_data[90207:90176] - in_data[90239:90208];
  assign out_data[45151:45120] = in_data[90271:90240] - in_data[90303:90272];
  assign out_data[45183:45152] = in_data[90335:90304] - in_data[90367:90336];
  assign out_data[45215:45184] = in_data[90399:90368] - in_data[90431:90400];
  assign out_data[45247:45216] = in_data[90463:90432] - in_data[90495:90464];
  assign out_data[45279:45248] = in_data[90527:90496] - in_data[90559:90528];
  assign out_data[45311:45280] = in_data[90591:90560] - in_data[90623:90592];
  assign out_data[45343:45312] = in_data[90655:90624] - in_data[90687:90656];
  assign out_data[45375:45344] = in_data[90719:90688] - in_data[90751:90720];
  assign out_data[45407:45376] = in_data[90783:90752] - in_data[90815:90784];
  assign out_data[4543:4512] = in_data[9055:9024] - in_data[9087:9056];
  assign out_data[45439:45408] = in_data[90847:90816] - in_data[90879:90848];
  assign out_data[45471:45440] = in_data[90911:90880] - in_data[90943:90912];
  assign out_data[45503:45472] = in_data[90975:90944] - in_data[91007:90976];
  assign out_data[45535:45504] = in_data[91039:91008] - in_data[91071:91040];
  assign out_data[45567:45536] = in_data[91103:91072] - in_data[91135:91104];
  assign out_data[45599:45568] = in_data[91167:91136] - in_data[91199:91168];
  assign out_data[45631:45600] = in_data[91231:91200] - in_data[91263:91232];
  assign out_data[45663:45632] = in_data[91295:91264] - in_data[91327:91296];
  assign out_data[45695:45664] = in_data[91359:91328] - in_data[91391:91360];
  assign out_data[45727:45696] = in_data[91423:91392] - in_data[91455:91424];
  assign out_data[4575:4544] = in_data[9119:9088] - in_data[9151:9120];
  assign out_data[45759:45728] = in_data[91487:91456] - in_data[91519:91488];
  assign out_data[45791:45760] = in_data[91551:91520] - in_data[91583:91552];
  assign out_data[45823:45792] = in_data[91615:91584] - in_data[91647:91616];
  assign out_data[45855:45824] = in_data[91679:91648] - in_data[91711:91680];
  assign out_data[45887:45856] = in_data[91743:91712] - in_data[91775:91744];
  assign out_data[45919:45888] = in_data[91807:91776] - in_data[91839:91808];
  assign out_data[45951:45920] = in_data[91871:91840] - in_data[91903:91872];
  assign out_data[45983:45952] = in_data[91935:91904] - in_data[91967:91936];
  assign out_data[46015:45984] = in_data[91999:91968] - in_data[92031:92000];
  assign out_data[46047:46016] = in_data[92063:92032] - in_data[92095:92064];
  assign out_data[4607:4576] = in_data[9183:9152] - in_data[9215:9184];
  assign out_data[46079:46048] = in_data[92127:92096] - in_data[92159:92128];
  assign out_data[46111:46080] = in_data[92191:92160] - in_data[92223:92192];
  assign out_data[46143:46112] = in_data[92255:92224] - in_data[92287:92256];
  assign out_data[46175:46144] = in_data[92319:92288] - in_data[92351:92320];
  assign out_data[46207:46176] = in_data[92383:92352] - in_data[92415:92384];
  assign out_data[46239:46208] = in_data[92447:92416] - in_data[92479:92448];
  assign out_data[46271:46240] = in_data[92511:92480] - in_data[92543:92512];
  assign out_data[46303:46272] = in_data[92575:92544] - in_data[92607:92576];
  assign out_data[46335:46304] = in_data[92639:92608] - in_data[92671:92640];
  assign out_data[46367:46336] = in_data[92703:92672] - in_data[92735:92704];
  assign out_data[4639:4608] = in_data[9247:9216] - in_data[9279:9248];
  assign out_data[46399:46368] = in_data[92767:92736] - in_data[92799:92768];
  assign out_data[46431:46400] = in_data[92831:92800] - in_data[92863:92832];
  assign out_data[46463:46432] = in_data[92895:92864] - in_data[92927:92896];
  assign out_data[46495:46464] = in_data[92959:92928] - in_data[92991:92960];
  assign out_data[46527:46496] = in_data[93023:92992] - in_data[93055:93024];
  assign out_data[46559:46528] = in_data[93087:93056] - in_data[93119:93088];
  assign out_data[46591:46560] = in_data[93151:93120] - in_data[93183:93152];
  assign out_data[46623:46592] = in_data[93215:93184] - in_data[93247:93216];
  assign out_data[46655:46624] = in_data[93279:93248] - in_data[93311:93280];
  assign out_data[46687:46656] = in_data[93343:93312] - in_data[93375:93344];
  assign out_data[4671:4640] = in_data[9311:9280] - in_data[9343:9312];
  assign out_data[46719:46688] = in_data[93407:93376] - in_data[93439:93408];
  assign out_data[46751:46720] = in_data[93471:93440] - in_data[93503:93472];
  assign out_data[46783:46752] = in_data[93535:93504] - in_data[93567:93536];
  assign out_data[46815:46784] = in_data[93599:93568] - in_data[93631:93600];
  assign out_data[46847:46816] = in_data[93663:93632] - in_data[93695:93664];
  assign out_data[46879:46848] = in_data[93727:93696] - in_data[93759:93728];
  assign out_data[46911:46880] = in_data[93791:93760] - in_data[93823:93792];
  assign out_data[46943:46912] = in_data[93855:93824] - in_data[93887:93856];
  assign out_data[46975:46944] = in_data[93919:93888] - in_data[93951:93920];
  assign out_data[47007:46976] = in_data[93983:93952] - in_data[94015:93984];
  assign out_data[4703:4672] = in_data[9375:9344] - in_data[9407:9376];
  assign out_data[47039:47008] = in_data[94047:94016] - in_data[94079:94048];
  assign out_data[47071:47040] = in_data[94111:94080] - in_data[94143:94112];
  assign out_data[47103:47072] = in_data[94175:94144] - in_data[94207:94176];
  assign out_data[47135:47104] = in_data[94239:94208] - in_data[94271:94240];
  assign out_data[47167:47136] = in_data[94303:94272] - in_data[94335:94304];
  assign out_data[47199:47168] = in_data[94367:94336] - in_data[94399:94368];
  assign out_data[47231:47200] = in_data[94431:94400] - in_data[94463:94432];
  assign out_data[47263:47232] = in_data[94495:94464] - in_data[94527:94496];
  assign out_data[47295:47264] = in_data[94559:94528] - in_data[94591:94560];
  assign out_data[47327:47296] = in_data[94623:94592] - in_data[94655:94624];
  assign out_data[4735:4704] = in_data[9439:9408] - in_data[9471:9440];
  assign out_data[47359:47328] = in_data[94687:94656] - in_data[94719:94688];
  assign out_data[47391:47360] = in_data[94751:94720] - in_data[94783:94752];
  assign out_data[47423:47392] = in_data[94815:94784] - in_data[94847:94816];
  assign out_data[47455:47424] = in_data[94879:94848] - in_data[94911:94880];
  assign out_data[47487:47456] = in_data[94943:94912] - in_data[94975:94944];
  assign out_data[47519:47488] = in_data[95007:94976] - in_data[95039:95008];
  assign out_data[47551:47520] = in_data[95071:95040] - in_data[95103:95072];
  assign out_data[47583:47552] = in_data[95135:95104] - in_data[95167:95136];
  assign out_data[47615:47584] = in_data[95199:95168] - in_data[95231:95200];
  assign out_data[47647:47616] = in_data[95263:95232] - in_data[95295:95264];
  assign out_data[4767:4736] = in_data[9503:9472] - in_data[9535:9504];
  assign out_data[47679:47648] = in_data[95327:95296] - in_data[95359:95328];
  assign out_data[47711:47680] = in_data[95391:95360] - in_data[95423:95392];
  assign out_data[47743:47712] = in_data[95455:95424] - in_data[95487:95456];
  assign out_data[47775:47744] = in_data[95519:95488] - in_data[95551:95520];
  assign out_data[47807:47776] = in_data[95583:95552] - in_data[95615:95584];
  assign out_data[47839:47808] = in_data[95647:95616] - in_data[95679:95648];
  assign out_data[47871:47840] = in_data[95711:95680] - in_data[95743:95712];
  assign out_data[47903:47872] = in_data[95775:95744] - in_data[95807:95776];
  assign out_data[47935:47904] = in_data[95839:95808] - in_data[95871:95840];
  assign out_data[47967:47936] = in_data[95903:95872] - in_data[95935:95904];
  assign out_data[479:448] = in_data[927:896] - in_data[959:928];
  assign out_data[4799:4768] = in_data[9567:9536] - in_data[9599:9568];
  assign out_data[47999:47968] = in_data[95967:95936] - in_data[95999:95968];
  assign out_data[48031:48000] = in_data[96031:96000] - in_data[96063:96032];
  assign out_data[48063:48032] = in_data[96095:96064] - in_data[96127:96096];
  assign out_data[48095:48064] = in_data[96159:96128] - in_data[96191:96160];
  assign out_data[48127:48096] = in_data[96223:96192] - in_data[96255:96224];
  assign out_data[48159:48128] = in_data[96287:96256] - in_data[96319:96288];
  assign out_data[48191:48160] = in_data[96351:96320] - in_data[96383:96352];
  assign out_data[48223:48192] = in_data[96415:96384] - in_data[96447:96416];
  assign out_data[48255:48224] = in_data[96479:96448] - in_data[96511:96480];
  assign out_data[48287:48256] = in_data[96543:96512] - in_data[96575:96544];
  assign out_data[4831:4800] = in_data[9631:9600] - in_data[9663:9632];
  assign out_data[48319:48288] = in_data[96607:96576] - in_data[96639:96608];
  assign out_data[48351:48320] = in_data[96671:96640] - in_data[96703:96672];
  assign out_data[48383:48352] = in_data[96735:96704] - in_data[96767:96736];
  assign out_data[48415:48384] = in_data[96799:96768] - in_data[96831:96800];
  assign out_data[48447:48416] = in_data[96863:96832] - in_data[96895:96864];
  assign out_data[48479:48448] = in_data[96927:96896] - in_data[96959:96928];
  assign out_data[48511:48480] = in_data[96991:96960] - in_data[97023:96992];
  assign out_data[48543:48512] = in_data[97055:97024] - in_data[97087:97056];
  assign out_data[48575:48544] = in_data[97119:97088] - in_data[97151:97120];
  assign out_data[48607:48576] = in_data[97183:97152] - in_data[97215:97184];
  assign out_data[4863:4832] = in_data[9695:9664] - in_data[9727:9696];
  assign out_data[48639:48608] = in_data[97247:97216] - in_data[97279:97248];
  assign out_data[48671:48640] = in_data[97311:97280] - in_data[97343:97312];
  assign out_data[48703:48672] = in_data[97375:97344] - in_data[97407:97376];
  assign out_data[48735:48704] = in_data[97439:97408] - in_data[97471:97440];
  assign out_data[48767:48736] = in_data[97503:97472] - in_data[97535:97504];
  assign out_data[48799:48768] = in_data[97567:97536] - in_data[97599:97568];
  assign out_data[48831:48800] = in_data[97631:97600] - in_data[97663:97632];
  assign out_data[48863:48832] = in_data[97695:97664] - in_data[97727:97696];
  assign out_data[48895:48864] = in_data[97759:97728] - in_data[97791:97760];
  assign out_data[48927:48896] = in_data[97823:97792] - in_data[97855:97824];
  assign out_data[4895:4864] = in_data[9759:9728] - in_data[9791:9760];
  assign out_data[48959:48928] = in_data[97887:97856] - in_data[97919:97888];
  assign out_data[48991:48960] = in_data[97951:97920] - in_data[97983:97952];
  assign out_data[49023:48992] = in_data[98015:97984] - in_data[98047:98016];
  assign out_data[49055:49024] = in_data[98079:98048] - in_data[98111:98080];
  assign out_data[49087:49056] = in_data[98143:98112] - in_data[98175:98144];
  assign out_data[49119:49088] = in_data[98207:98176] - in_data[98239:98208];
  assign out_data[49151:49120] = in_data[98271:98240] - in_data[98303:98272];
  assign out_data[49183:49152] = in_data[98335:98304] - in_data[98367:98336];
  assign out_data[49215:49184] = in_data[98399:98368] - in_data[98431:98400];
  assign out_data[49247:49216] = in_data[98463:98432] - in_data[98495:98464];
  assign out_data[4927:4896] = in_data[9823:9792] - in_data[9855:9824];
  assign out_data[49279:49248] = in_data[98527:98496] - in_data[98559:98528];
  assign out_data[49311:49280] = in_data[98591:98560] - in_data[98623:98592];
  assign out_data[49343:49312] = in_data[98655:98624] - in_data[98687:98656];
  assign out_data[49375:49344] = in_data[98719:98688] - in_data[98751:98720];
  assign out_data[49407:49376] = in_data[98783:98752] - in_data[98815:98784];
  assign out_data[49439:49408] = in_data[98847:98816] - in_data[98879:98848];
  assign out_data[49471:49440] = in_data[98911:98880] - in_data[98943:98912];
  assign out_data[49503:49472] = in_data[98975:98944] - in_data[99007:98976];
  assign out_data[49535:49504] = in_data[99039:99008] - in_data[99071:99040];
  assign out_data[49567:49536] = in_data[99103:99072] - in_data[99135:99104];
  assign out_data[4959:4928] = in_data[9887:9856] - in_data[9919:9888];
  assign out_data[49599:49568] = in_data[99167:99136] - in_data[99199:99168];
  assign out_data[49631:49600] = in_data[99231:99200] - in_data[99263:99232];
  assign out_data[49663:49632] = in_data[99295:99264] - in_data[99327:99296];
  assign out_data[49695:49664] = in_data[99359:99328] - in_data[99391:99360];
  assign out_data[49727:49696] = in_data[99423:99392] - in_data[99455:99424];
  assign out_data[49759:49728] = in_data[99487:99456] - in_data[99519:99488];
  assign out_data[49791:49760] = in_data[99551:99520] - in_data[99583:99552];
  assign out_data[49823:49792] = in_data[99615:99584] - in_data[99647:99616];
  assign out_data[49855:49824] = in_data[99679:99648] - in_data[99711:99680];
  assign out_data[49887:49856] = in_data[99743:99712] - in_data[99775:99744];
  assign out_data[4991:4960] = in_data[9951:9920] - in_data[9983:9952];
  assign out_data[49919:49888] = in_data[99807:99776] - in_data[99839:99808];
  assign out_data[49951:49920] = in_data[99871:99840] - in_data[99903:99872];
  assign out_data[49983:49952] = in_data[99935:99904] - in_data[99967:99936];
  assign out_data[50015:49984] = in_data[99999:99968] - in_data[100031:100000];
  assign out_data[50047:50016] = in_data[100063:100032] - in_data[100095:100064];
  assign out_data[50079:50048] = in_data[100127:100096] - in_data[100159:100128];
  assign out_data[50111:50080] = in_data[100191:100160] - in_data[100223:100192];
  assign out_data[50143:50112] = in_data[100255:100224] - in_data[100287:100256];
  assign out_data[50175:50144] = in_data[100319:100288] - in_data[100351:100320];
  assign out_data[50207:50176] = in_data[100383:100352] - in_data[100415:100384];
  assign out_data[5023:4992] = in_data[10015:9984] - in_data[10047:10016];
  assign out_data[50239:50208] = in_data[100447:100416] - in_data[100479:100448];
  assign out_data[50271:50240] = in_data[100511:100480] - in_data[100543:100512];
  assign out_data[50303:50272] = in_data[100575:100544] - in_data[100607:100576];
  assign out_data[50335:50304] = in_data[100639:100608] - in_data[100671:100640];
  assign out_data[50367:50336] = in_data[100703:100672] - in_data[100735:100704];
  assign out_data[50399:50368] = in_data[100767:100736] - in_data[100799:100768];
  assign out_data[50431:50400] = in_data[100831:100800] - in_data[100863:100832];
  assign out_data[50463:50432] = in_data[100895:100864] - in_data[100927:100896];
  assign out_data[50495:50464] = in_data[100959:100928] - in_data[100991:100960];
  assign out_data[50527:50496] = in_data[101023:100992] - in_data[101055:101024];
  assign out_data[5055:5024] = in_data[10079:10048] - in_data[10111:10080];
  assign out_data[50559:50528] = in_data[101087:101056] - in_data[101119:101088];
  assign out_data[50591:50560] = in_data[101151:101120] - in_data[101183:101152];
  assign out_data[50623:50592] = in_data[101215:101184] - in_data[101247:101216];
  assign out_data[50655:50624] = in_data[101279:101248] - in_data[101311:101280];
  assign out_data[50687:50656] = in_data[101343:101312] - in_data[101375:101344];
  assign out_data[50719:50688] = in_data[101407:101376] - in_data[101439:101408];
  assign out_data[50751:50720] = in_data[101471:101440] - in_data[101503:101472];
  assign out_data[50783:50752] = in_data[101535:101504] - in_data[101567:101536];
  assign out_data[50815:50784] = in_data[101599:101568] - in_data[101631:101600];
  assign out_data[50847:50816] = in_data[101663:101632] - in_data[101695:101664];
  assign out_data[5087:5056] = in_data[10143:10112] - in_data[10175:10144];
  assign out_data[50879:50848] = in_data[101727:101696] - in_data[101759:101728];
  assign out_data[50911:50880] = in_data[101791:101760] - in_data[101823:101792];
  assign out_data[50943:50912] = in_data[101855:101824] - in_data[101887:101856];
  assign out_data[50975:50944] = in_data[101919:101888] - in_data[101951:101920];
  assign out_data[51007:50976] = in_data[101983:101952] - in_data[102015:101984];
  assign out_data[51039:51008] = in_data[102047:102016] - in_data[102079:102048];
  assign out_data[51071:51040] = in_data[102111:102080] - in_data[102143:102112];
  assign out_data[51103:51072] = in_data[102175:102144] - in_data[102207:102176];
  assign out_data[51135:51104] = in_data[102239:102208] - in_data[102271:102240];
  assign out_data[51167:51136] = in_data[102303:102272] - in_data[102335:102304];
  assign out_data[511:480] = in_data[991:960] - in_data[1023:992];
  assign out_data[5119:5088] = in_data[10207:10176] - in_data[10239:10208];
  assign out_data[51199:51168] = in_data[102367:102336] - in_data[102399:102368];
  assign out_data[51231:51200] = in_data[102431:102400] - in_data[102463:102432];
  assign out_data[51263:51232] = in_data[102495:102464] - in_data[102527:102496];
  assign out_data[51295:51264] = in_data[102559:102528] - in_data[102591:102560];
  assign out_data[51327:51296] = in_data[102623:102592] - in_data[102655:102624];
  assign out_data[51359:51328] = in_data[102687:102656] - in_data[102719:102688];
  assign out_data[51391:51360] = in_data[102751:102720] - in_data[102783:102752];
  assign out_data[51423:51392] = in_data[102815:102784] - in_data[102847:102816];
  assign out_data[51455:51424] = in_data[102879:102848] - in_data[102911:102880];
  assign out_data[51487:51456] = in_data[102943:102912] - in_data[102975:102944];
  assign out_data[5151:5120] = in_data[10271:10240] - in_data[10303:10272];
  assign out_data[51519:51488] = in_data[103007:102976] - in_data[103039:103008];
  assign out_data[51551:51520] = in_data[103071:103040] - in_data[103103:103072];
  assign out_data[51583:51552] = in_data[103135:103104] - in_data[103167:103136];
  assign out_data[51615:51584] = in_data[103199:103168] - in_data[103231:103200];
  assign out_data[51647:51616] = in_data[103263:103232] - in_data[103295:103264];
  assign out_data[51679:51648] = in_data[103327:103296] - in_data[103359:103328];
  assign out_data[51711:51680] = in_data[103391:103360] - in_data[103423:103392];
  assign out_data[51743:51712] = in_data[103455:103424] - in_data[103487:103456];
  assign out_data[51775:51744] = in_data[103519:103488] - in_data[103551:103520];
  assign out_data[51807:51776] = in_data[103583:103552] - in_data[103615:103584];
  assign out_data[5183:5152] = in_data[10335:10304] - in_data[10367:10336];
  assign out_data[51839:51808] = in_data[103647:103616] - in_data[103679:103648];
  assign out_data[51871:51840] = in_data[103711:103680] - in_data[103743:103712];
  assign out_data[51903:51872] = in_data[103775:103744] - in_data[103807:103776];
  assign out_data[51935:51904] = in_data[103839:103808] - in_data[103871:103840];
  assign out_data[51967:51936] = in_data[103903:103872] - in_data[103935:103904];
  assign out_data[51999:51968] = in_data[103967:103936] - in_data[103999:103968];
  assign out_data[52031:52000] = in_data[104031:104000] - in_data[104063:104032];
  assign out_data[52063:52032] = in_data[104095:104064] - in_data[104127:104096];
  assign out_data[52095:52064] = in_data[104159:104128] - in_data[104191:104160];
  assign out_data[52127:52096] = in_data[104223:104192] - in_data[104255:104224];
  assign out_data[5215:5184] = in_data[10399:10368] - in_data[10431:10400];
  assign out_data[52159:52128] = in_data[104287:104256] - in_data[104319:104288];
  assign out_data[52191:52160] = in_data[104351:104320] - in_data[104383:104352];
  assign out_data[52223:52192] = in_data[104415:104384] - in_data[104447:104416];
  assign out_data[52255:52224] = in_data[104479:104448] - in_data[104511:104480];
  assign out_data[52287:52256] = in_data[104543:104512] - in_data[104575:104544];
  assign out_data[52319:52288] = in_data[104607:104576] - in_data[104639:104608];
  assign out_data[52351:52320] = in_data[104671:104640] - in_data[104703:104672];
  assign out_data[52383:52352] = in_data[104735:104704] - in_data[104767:104736];
  assign out_data[52415:52384] = in_data[104799:104768] - in_data[104831:104800];
  assign out_data[52447:52416] = in_data[104863:104832] - in_data[104895:104864];
  assign out_data[5247:5216] = in_data[10463:10432] - in_data[10495:10464];
  assign out_data[52479:52448] = in_data[104927:104896] - in_data[104959:104928];
  assign out_data[52511:52480] = in_data[104991:104960] - in_data[105023:104992];
  assign out_data[52543:52512] = in_data[105055:105024] - in_data[105087:105056];
  assign out_data[52575:52544] = in_data[105119:105088] - in_data[105151:105120];
  assign out_data[52607:52576] = in_data[105183:105152] - in_data[105215:105184];
  assign out_data[52639:52608] = in_data[105247:105216] - in_data[105279:105248];
  assign out_data[52671:52640] = in_data[105311:105280] - in_data[105343:105312];
  assign out_data[52703:52672] = in_data[105375:105344] - in_data[105407:105376];
  assign out_data[52735:52704] = in_data[105439:105408] - in_data[105471:105440];
  assign out_data[52767:52736] = in_data[105503:105472] - in_data[105535:105504];
  assign out_data[5279:5248] = in_data[10527:10496] - in_data[10559:10528];
  assign out_data[52799:52768] = in_data[105567:105536] - in_data[105599:105568];
  assign out_data[52831:52800] = in_data[105631:105600] - in_data[105663:105632];
  assign out_data[52863:52832] = in_data[105695:105664] - in_data[105727:105696];
  assign out_data[52895:52864] = in_data[105759:105728] - in_data[105791:105760];
  assign out_data[52927:52896] = in_data[105823:105792] - in_data[105855:105824];
  assign out_data[52959:52928] = in_data[105887:105856] - in_data[105919:105888];
  assign out_data[52991:52960] = in_data[105951:105920] - in_data[105983:105952];
  assign out_data[53023:52992] = in_data[106015:105984] - in_data[106047:106016];
  assign out_data[53055:53024] = in_data[106079:106048] - in_data[106111:106080];
  assign out_data[53087:53056] = in_data[106143:106112] - in_data[106175:106144];
  assign out_data[5311:5280] = in_data[10591:10560] - in_data[10623:10592];
  assign out_data[53119:53088] = in_data[106207:106176] - in_data[106239:106208];
  assign out_data[53151:53120] = in_data[106271:106240] - in_data[106303:106272];
  assign out_data[53183:53152] = in_data[106335:106304] - in_data[106367:106336];
  assign out_data[53215:53184] = in_data[106399:106368] - in_data[106431:106400];
  assign out_data[53247:53216] = in_data[106463:106432] - in_data[106495:106464];
  assign out_data[53279:53248] = in_data[106527:106496] - in_data[106559:106528];
  assign out_data[53311:53280] = in_data[106591:106560] - in_data[106623:106592];
  assign out_data[53343:53312] = in_data[106655:106624] - in_data[106687:106656];
  assign out_data[53375:53344] = in_data[106719:106688] - in_data[106751:106720];
  assign out_data[53407:53376] = in_data[106783:106752] - in_data[106815:106784];
  assign out_data[5343:5312] = in_data[10655:10624] - in_data[10687:10656];
  assign out_data[53439:53408] = in_data[106847:106816] - in_data[106879:106848];
  assign out_data[53471:53440] = in_data[106911:106880] - in_data[106943:106912];
  assign out_data[53503:53472] = in_data[106975:106944] - in_data[107007:106976];
  assign out_data[53535:53504] = in_data[107039:107008] - in_data[107071:107040];
  assign out_data[53567:53536] = in_data[107103:107072] - in_data[107135:107104];
  assign out_data[53599:53568] = in_data[107167:107136] - in_data[107199:107168];
  assign out_data[53631:53600] = in_data[107231:107200] - in_data[107263:107232];
  assign out_data[53663:53632] = in_data[107295:107264] - in_data[107327:107296];
  assign out_data[53695:53664] = in_data[107359:107328] - in_data[107391:107360];
  assign out_data[53727:53696] = in_data[107423:107392] - in_data[107455:107424];
  assign out_data[5375:5344] = in_data[10719:10688] - in_data[10751:10720];
  assign out_data[53759:53728] = in_data[107487:107456] - in_data[107519:107488];
  assign out_data[53791:53760] = in_data[107551:107520] - in_data[107583:107552];
  assign out_data[53823:53792] = in_data[107615:107584] - in_data[107647:107616];
  assign out_data[53855:53824] = in_data[107679:107648] - in_data[107711:107680];
  assign out_data[53887:53856] = in_data[107743:107712] - in_data[107775:107744];
  assign out_data[53919:53888] = in_data[107807:107776] - in_data[107839:107808];
  assign out_data[53951:53920] = in_data[107871:107840] - in_data[107903:107872];
  assign out_data[53983:53952] = in_data[107935:107904] - in_data[107967:107936];
  assign out_data[54015:53984] = in_data[107999:107968] - in_data[108031:108000];
  assign out_data[54047:54016] = in_data[108063:108032] - in_data[108095:108064];
  assign out_data[5407:5376] = in_data[10783:10752] - in_data[10815:10784];
  assign out_data[54079:54048] = in_data[108127:108096] - in_data[108159:108128];
  assign out_data[54111:54080] = in_data[108191:108160] - in_data[108223:108192];
  assign out_data[54143:54112] = in_data[108255:108224] - in_data[108287:108256];
  assign out_data[54175:54144] = in_data[108319:108288] - in_data[108351:108320];
  assign out_data[54207:54176] = in_data[108383:108352] - in_data[108415:108384];
  assign out_data[54239:54208] = in_data[108447:108416] - in_data[108479:108448];
  assign out_data[54271:54240] = in_data[108511:108480] - in_data[108543:108512];
  assign out_data[54303:54272] = in_data[108575:108544] - in_data[108607:108576];
  assign out_data[54335:54304] = in_data[108639:108608] - in_data[108671:108640];
  assign out_data[54367:54336] = in_data[108703:108672] - in_data[108735:108704];
  assign out_data[543:512] = in_data[1055:1024] - in_data[1087:1056];
  assign out_data[5439:5408] = in_data[10847:10816] - in_data[10879:10848];
  assign out_data[54399:54368] = in_data[108767:108736] - in_data[108799:108768];
  assign out_data[54431:54400] = in_data[108831:108800] - in_data[108863:108832];
  assign out_data[54463:54432] = in_data[108895:108864] - in_data[108927:108896];
  assign out_data[54495:54464] = in_data[108959:108928] - in_data[108991:108960];
  assign out_data[54527:54496] = in_data[109023:108992] - in_data[109055:109024];
  assign out_data[54559:54528] = in_data[109087:109056] - in_data[109119:109088];
  assign out_data[54591:54560] = in_data[109151:109120] - in_data[109183:109152];
  assign out_data[54623:54592] = in_data[109215:109184] - in_data[109247:109216];
  assign out_data[54655:54624] = in_data[109279:109248] - in_data[109311:109280];
  assign out_data[54687:54656] = in_data[109343:109312] - in_data[109375:109344];
  assign out_data[5471:5440] = in_data[10911:10880] - in_data[10943:10912];
  assign out_data[54719:54688] = in_data[109407:109376] - in_data[109439:109408];
  assign out_data[54751:54720] = in_data[109471:109440] - in_data[109503:109472];
  assign out_data[54783:54752] = in_data[109535:109504] - in_data[109567:109536];
  assign out_data[54815:54784] = in_data[109599:109568] - in_data[109631:109600];
  assign out_data[54847:54816] = in_data[109663:109632] - in_data[109695:109664];
  assign out_data[54879:54848] = in_data[109727:109696] - in_data[109759:109728];
  assign out_data[54911:54880] = in_data[109791:109760] - in_data[109823:109792];
  assign out_data[54943:54912] = in_data[109855:109824] - in_data[109887:109856];
  assign out_data[54975:54944] = in_data[109919:109888] - in_data[109951:109920];
  assign out_data[55007:54976] = in_data[109983:109952] - in_data[110015:109984];
  assign out_data[5503:5472] = in_data[10975:10944] - in_data[11007:10976];
  assign out_data[55039:55008] = in_data[110047:110016] - in_data[110079:110048];
  assign out_data[55071:55040] = in_data[110111:110080] - in_data[110143:110112];
  assign out_data[55103:55072] = in_data[110175:110144] - in_data[110207:110176];
  assign out_data[55135:55104] = in_data[110239:110208] - in_data[110271:110240];
  assign out_data[55167:55136] = in_data[110303:110272] - in_data[110335:110304];
  assign out_data[55199:55168] = in_data[110367:110336] - in_data[110399:110368];
  assign out_data[55231:55200] = in_data[110431:110400] - in_data[110463:110432];
  assign out_data[55263:55232] = in_data[110495:110464] - in_data[110527:110496];
  assign out_data[55295:55264] = in_data[110559:110528] - in_data[110591:110560];
  assign out_data[55327:55296] = in_data[110623:110592] - in_data[110655:110624];
  assign out_data[5535:5504] = in_data[11039:11008] - in_data[11071:11040];
  assign out_data[55359:55328] = in_data[110687:110656] - in_data[110719:110688];
  assign out_data[55391:55360] = in_data[110751:110720] - in_data[110783:110752];
  assign out_data[55423:55392] = in_data[110815:110784] - in_data[110847:110816];
  assign out_data[55455:55424] = in_data[110879:110848] - in_data[110911:110880];
  assign out_data[55487:55456] = in_data[110943:110912] - in_data[110975:110944];
  assign out_data[55519:55488] = in_data[111007:110976] - in_data[111039:111008];
  assign out_data[55551:55520] = in_data[111071:111040] - in_data[111103:111072];
  assign out_data[55583:55552] = in_data[111135:111104] - in_data[111167:111136];
  assign out_data[55615:55584] = in_data[111199:111168] - in_data[111231:111200];
  assign out_data[55647:55616] = in_data[111263:111232] - in_data[111295:111264];
  assign out_data[5567:5536] = in_data[11103:11072] - in_data[11135:11104];
  assign out_data[55679:55648] = in_data[111327:111296] - in_data[111359:111328];
  assign out_data[55711:55680] = in_data[111391:111360] - in_data[111423:111392];
  assign out_data[55743:55712] = in_data[111455:111424] - in_data[111487:111456];
  assign out_data[55775:55744] = in_data[111519:111488] - in_data[111551:111520];
  assign out_data[55807:55776] = in_data[111583:111552] - in_data[111615:111584];
  assign out_data[55839:55808] = in_data[111647:111616] - in_data[111679:111648];
  assign out_data[55871:55840] = in_data[111711:111680] - in_data[111743:111712];
  assign out_data[55903:55872] = in_data[111775:111744] - in_data[111807:111776];
  assign out_data[55935:55904] = in_data[111839:111808] - in_data[111871:111840];
  assign out_data[55967:55936] = in_data[111903:111872] - in_data[111935:111904];
  assign out_data[5599:5568] = in_data[11167:11136] - in_data[11199:11168];
  assign out_data[55999:55968] = in_data[111967:111936] - in_data[111999:111968];
  assign out_data[56031:56000] = in_data[112031:112000] - in_data[112063:112032];
  assign out_data[56063:56032] = in_data[112095:112064] - in_data[112127:112096];
  assign out_data[56095:56064] = in_data[112159:112128] - in_data[112191:112160];
  assign out_data[56127:56096] = in_data[112223:112192] - in_data[112255:112224];
  assign out_data[56159:56128] = in_data[112287:112256] - in_data[112319:112288];
  assign out_data[56191:56160] = in_data[112351:112320] - in_data[112383:112352];
  assign out_data[56223:56192] = in_data[112415:112384] - in_data[112447:112416];
  assign out_data[56255:56224] = in_data[112479:112448] - in_data[112511:112480];
  assign out_data[56287:56256] = in_data[112543:112512] - in_data[112575:112544];
  assign out_data[5631:5600] = in_data[11231:11200] - in_data[11263:11232];
  assign out_data[56319:56288] = in_data[112607:112576] - in_data[112639:112608];
  assign out_data[56351:56320] = in_data[112671:112640] - in_data[112703:112672];
  assign out_data[56383:56352] = in_data[112735:112704] - in_data[112767:112736];
  assign out_data[56415:56384] = in_data[112799:112768] - in_data[112831:112800];
  assign out_data[56447:56416] = in_data[112863:112832] - in_data[112895:112864];
  assign out_data[56479:56448] = in_data[112927:112896] - in_data[112959:112928];
  assign out_data[56511:56480] = in_data[112991:112960] - in_data[113023:112992];
  assign out_data[56543:56512] = in_data[113055:113024] - in_data[113087:113056];
  assign out_data[56575:56544] = in_data[113119:113088] - in_data[113151:113120];
  assign out_data[56607:56576] = in_data[113183:113152] - in_data[113215:113184];
  assign out_data[5663:5632] = in_data[11295:11264] - in_data[11327:11296];
  assign out_data[56639:56608] = in_data[113247:113216] - in_data[113279:113248];
  assign out_data[56671:56640] = in_data[113311:113280] - in_data[113343:113312];
  assign out_data[56703:56672] = in_data[113375:113344] - in_data[113407:113376];
  assign out_data[56735:56704] = in_data[113439:113408] - in_data[113471:113440];
  assign out_data[56767:56736] = in_data[113503:113472] - in_data[113535:113504];
  assign out_data[56799:56768] = in_data[113567:113536] - in_data[113599:113568];
  assign out_data[56831:56800] = in_data[113631:113600] - in_data[113663:113632];
  assign out_data[56863:56832] = in_data[113695:113664] - in_data[113727:113696];
  assign out_data[56895:56864] = in_data[113759:113728] - in_data[113791:113760];
  assign out_data[56927:56896] = in_data[113823:113792] - in_data[113855:113824];
  assign out_data[5695:5664] = in_data[11359:11328] - in_data[11391:11360];
  assign out_data[56959:56928] = in_data[113887:113856] - in_data[113919:113888];
  assign out_data[56991:56960] = in_data[113951:113920] - in_data[113983:113952];
  assign out_data[57023:56992] = in_data[114015:113984] - in_data[114047:114016];
  assign out_data[57055:57024] = in_data[114079:114048] - in_data[114111:114080];
  assign out_data[57087:57056] = in_data[114143:114112] - in_data[114175:114144];
  assign out_data[57119:57088] = in_data[114207:114176] - in_data[114239:114208];
  assign out_data[57151:57120] = in_data[114271:114240] - in_data[114303:114272];
  assign out_data[57183:57152] = in_data[114335:114304] - in_data[114367:114336];
  assign out_data[57215:57184] = in_data[114399:114368] - in_data[114431:114400];
  assign out_data[57247:57216] = in_data[114463:114432] - in_data[114495:114464];
  assign out_data[5727:5696] = in_data[11423:11392] - in_data[11455:11424];
  assign out_data[57279:57248] = in_data[114527:114496] - in_data[114559:114528];
  assign out_data[57311:57280] = in_data[114591:114560] - in_data[114623:114592];
  assign out_data[57343:57312] = in_data[114655:114624] - in_data[114687:114656];
  assign out_data[57375:57344] = in_data[114719:114688] - in_data[114751:114720];
  assign out_data[57407:57376] = in_data[114783:114752] - in_data[114815:114784];
  assign out_data[57439:57408] = in_data[114847:114816] - in_data[114879:114848];
  assign out_data[57471:57440] = in_data[114911:114880] - in_data[114943:114912];
  assign out_data[57503:57472] = in_data[114975:114944] - in_data[115007:114976];
  assign out_data[57535:57504] = in_data[115039:115008] - in_data[115071:115040];
  assign out_data[57567:57536] = in_data[115103:115072] - in_data[115135:115104];
  assign out_data[575:544] = in_data[1119:1088] - in_data[1151:1120];
  assign out_data[5759:5728] = in_data[11487:11456] - in_data[11519:11488];
  assign out_data[57599:57568] = in_data[115167:115136] - in_data[115199:115168];
  assign out_data[57631:57600] = in_data[115231:115200] - in_data[115263:115232];
  assign out_data[57663:57632] = in_data[115295:115264] - in_data[115327:115296];
  assign out_data[57695:57664] = in_data[115359:115328] - in_data[115391:115360];
  assign out_data[57727:57696] = in_data[115423:115392] - in_data[115455:115424];
  assign out_data[57759:57728] = in_data[115487:115456] - in_data[115519:115488];
  assign out_data[57791:57760] = in_data[115551:115520] - in_data[115583:115552];
  assign out_data[57823:57792] = in_data[115615:115584] - in_data[115647:115616];
  assign out_data[57855:57824] = in_data[115679:115648] - in_data[115711:115680];
  assign out_data[57887:57856] = in_data[115743:115712] - in_data[115775:115744];
  assign out_data[5791:5760] = in_data[11551:11520] - in_data[11583:11552];
  assign out_data[57919:57888] = in_data[115807:115776] - in_data[115839:115808];
  assign out_data[57951:57920] = in_data[115871:115840] - in_data[115903:115872];
  assign out_data[57983:57952] = in_data[115935:115904] - in_data[115967:115936];
  assign out_data[58015:57984] = in_data[115999:115968] - in_data[116031:116000];
  assign out_data[58047:58016] = in_data[116063:116032] - in_data[116095:116064];
  assign out_data[58079:58048] = in_data[116127:116096] - in_data[116159:116128];
  assign out_data[58111:58080] = in_data[116191:116160] - in_data[116223:116192];
  assign out_data[58143:58112] = in_data[116255:116224] - in_data[116287:116256];
  assign out_data[58175:58144] = in_data[116319:116288] - in_data[116351:116320];
  assign out_data[58207:58176] = in_data[116383:116352] - in_data[116415:116384];
  assign out_data[5823:5792] = in_data[11615:11584] - in_data[11647:11616];
  assign out_data[58239:58208] = in_data[116447:116416] - in_data[116479:116448];
  assign out_data[58271:58240] = in_data[116511:116480] - in_data[116543:116512];
  assign out_data[58303:58272] = in_data[116575:116544] - in_data[116607:116576];
  assign out_data[58335:58304] = in_data[116639:116608] - in_data[116671:116640];
  assign out_data[58367:58336] = in_data[116703:116672] - in_data[116735:116704];
  assign out_data[58399:58368] = in_data[116767:116736] - in_data[116799:116768];
  assign out_data[58431:58400] = in_data[116831:116800] - in_data[116863:116832];
  assign out_data[58463:58432] = in_data[116895:116864] - in_data[116927:116896];
  assign out_data[58495:58464] = in_data[116959:116928] - in_data[116991:116960];
  assign out_data[58527:58496] = in_data[117023:116992] - in_data[117055:117024];
  assign out_data[5855:5824] = in_data[11679:11648] - in_data[11711:11680];
  assign out_data[58559:58528] = in_data[117087:117056] - in_data[117119:117088];
  assign out_data[58591:58560] = in_data[117151:117120] - in_data[117183:117152];
  assign out_data[58623:58592] = in_data[117215:117184] - in_data[117247:117216];
  assign out_data[58655:58624] = in_data[117279:117248] - in_data[117311:117280];
  assign out_data[58687:58656] = in_data[117343:117312] - in_data[117375:117344];
  assign out_data[58719:58688] = in_data[117407:117376] - in_data[117439:117408];
  assign out_data[58751:58720] = in_data[117471:117440] - in_data[117503:117472];
  assign out_data[58783:58752] = in_data[117535:117504] - in_data[117567:117536];
  assign out_data[58815:58784] = in_data[117599:117568] - in_data[117631:117600];
  assign out_data[58847:58816] = in_data[117663:117632] - in_data[117695:117664];
  assign out_data[5887:5856] = in_data[11743:11712] - in_data[11775:11744];
  assign out_data[58879:58848] = in_data[117727:117696] - in_data[117759:117728];
  assign out_data[58911:58880] = in_data[117791:117760] - in_data[117823:117792];
  assign out_data[58943:58912] = in_data[117855:117824] - in_data[117887:117856];
  assign out_data[58975:58944] = in_data[117919:117888] - in_data[117951:117920];
  assign out_data[59007:58976] = in_data[117983:117952] - in_data[118015:117984];
  assign out_data[59039:59008] = in_data[118047:118016] - in_data[118079:118048];
  assign out_data[59071:59040] = in_data[118111:118080] - in_data[118143:118112];
  assign out_data[59103:59072] = in_data[118175:118144] - in_data[118207:118176];
  assign out_data[59135:59104] = in_data[118239:118208] - in_data[118271:118240];
  assign out_data[59167:59136] = in_data[118303:118272] - in_data[118335:118304];
  assign out_data[5919:5888] = in_data[11807:11776] - in_data[11839:11808];
  assign out_data[59199:59168] = in_data[118367:118336] - in_data[118399:118368];
  assign out_data[59231:59200] = in_data[118431:118400] - in_data[118463:118432];
  assign out_data[59263:59232] = in_data[118495:118464] - in_data[118527:118496];
  assign out_data[59295:59264] = in_data[118559:118528] - in_data[118591:118560];
  assign out_data[59327:59296] = in_data[118623:118592] - in_data[118655:118624];
  assign out_data[59359:59328] = in_data[118687:118656] - in_data[118719:118688];
  assign out_data[59391:59360] = in_data[118751:118720] - in_data[118783:118752];
  assign out_data[59423:59392] = in_data[118815:118784] - in_data[118847:118816];
  assign out_data[59455:59424] = in_data[118879:118848] - in_data[118911:118880];
  assign out_data[59487:59456] = in_data[118943:118912] - in_data[118975:118944];
  assign out_data[5951:5920] = in_data[11871:11840] - in_data[11903:11872];
  assign out_data[59519:59488] = in_data[119007:118976] - in_data[119039:119008];
  assign out_data[59551:59520] = in_data[119071:119040] - in_data[119103:119072];
  assign out_data[59583:59552] = in_data[119135:119104] - in_data[119167:119136];
  assign out_data[59615:59584] = in_data[119199:119168] - in_data[119231:119200];
  assign out_data[59647:59616] = in_data[119263:119232] - in_data[119295:119264];
  assign out_data[59679:59648] = in_data[119327:119296] - in_data[119359:119328];
  assign out_data[59711:59680] = in_data[119391:119360] - in_data[119423:119392];
  assign out_data[59743:59712] = in_data[119455:119424] - in_data[119487:119456];
  assign out_data[59775:59744] = in_data[119519:119488] - in_data[119551:119520];
  assign out_data[59807:59776] = in_data[119583:119552] - in_data[119615:119584];
  assign out_data[5983:5952] = in_data[11935:11904] - in_data[11967:11936];
  assign out_data[59839:59808] = in_data[119647:119616] - in_data[119679:119648];
  assign out_data[59871:59840] = in_data[119711:119680] - in_data[119743:119712];
  assign out_data[59903:59872] = in_data[119775:119744] - in_data[119807:119776];
  assign out_data[59935:59904] = in_data[119839:119808] - in_data[119871:119840];
  assign out_data[59967:59936] = in_data[119903:119872] - in_data[119935:119904];
  assign out_data[59999:59968] = in_data[119967:119936] - in_data[119999:119968];
  assign out_data[60031:60000] = in_data[120031:120000] - in_data[120063:120032];
  assign out_data[60063:60032] = in_data[120095:120064] - in_data[120127:120096];
  assign out_data[60095:60064] = in_data[120159:120128] - in_data[120191:120160];
  assign out_data[60127:60096] = in_data[120223:120192] - in_data[120255:120224];
  assign out_data[6015:5984] = in_data[11999:11968] - in_data[12031:12000];
  assign out_data[60159:60128] = in_data[120287:120256] - in_data[120319:120288];
  assign out_data[60191:60160] = in_data[120351:120320] - in_data[120383:120352];
  assign out_data[60223:60192] = in_data[120415:120384] - in_data[120447:120416];
  assign out_data[60255:60224] = in_data[120479:120448] - in_data[120511:120480];
  assign out_data[60287:60256] = in_data[120543:120512] - in_data[120575:120544];
  assign out_data[60319:60288] = in_data[120607:120576] - in_data[120639:120608];
  assign out_data[60351:60320] = in_data[120671:120640] - in_data[120703:120672];
  assign out_data[60383:60352] = in_data[120735:120704] - in_data[120767:120736];
  assign out_data[60415:60384] = in_data[120799:120768] - in_data[120831:120800];
  assign out_data[60447:60416] = in_data[120863:120832] - in_data[120895:120864];
  assign out_data[6047:6016] = in_data[12063:12032] - in_data[12095:12064];
  assign out_data[60479:60448] = in_data[120927:120896] - in_data[120959:120928];
  assign out_data[60511:60480] = in_data[120991:120960] - in_data[121023:120992];
  assign out_data[60543:60512] = in_data[121055:121024] - in_data[121087:121056];
  assign out_data[60575:60544] = in_data[121119:121088] - in_data[121151:121120];
  assign out_data[60607:60576] = in_data[121183:121152] - in_data[121215:121184];
  assign out_data[60639:60608] = in_data[121247:121216] - in_data[121279:121248];
  assign out_data[60671:60640] = in_data[121311:121280] - in_data[121343:121312];
  assign out_data[60703:60672] = in_data[121375:121344] - in_data[121407:121376];
  assign out_data[60735:60704] = in_data[121439:121408] - in_data[121471:121440];
  assign out_data[60767:60736] = in_data[121503:121472] - in_data[121535:121504];
  assign out_data[607:576] = in_data[1183:1152] - in_data[1215:1184];
  assign out_data[6079:6048] = in_data[12127:12096] - in_data[12159:12128];
  assign out_data[60799:60768] = in_data[121567:121536] - in_data[121599:121568];
  assign out_data[60831:60800] = in_data[121631:121600] - in_data[121663:121632];
  assign out_data[60863:60832] = in_data[121695:121664] - in_data[121727:121696];
  assign out_data[60895:60864] = in_data[121759:121728] - in_data[121791:121760];
  assign out_data[60927:60896] = in_data[121823:121792] - in_data[121855:121824];
  assign out_data[60959:60928] = in_data[121887:121856] - in_data[121919:121888];
  assign out_data[60991:60960] = in_data[121951:121920] - in_data[121983:121952];
  assign out_data[61023:60992] = in_data[122015:121984] - in_data[122047:122016];
  assign out_data[61055:61024] = in_data[122079:122048] - in_data[122111:122080];
  assign out_data[61087:61056] = in_data[122143:122112] - in_data[122175:122144];
  assign out_data[6111:6080] = in_data[12191:12160] - in_data[12223:12192];
  assign out_data[61119:61088] = in_data[122207:122176] - in_data[122239:122208];
  assign out_data[61151:61120] = in_data[122271:122240] - in_data[122303:122272];
  assign out_data[61183:61152] = in_data[122335:122304] - in_data[122367:122336];
  assign out_data[61215:61184] = in_data[122399:122368] - in_data[122431:122400];
  assign out_data[61247:61216] = in_data[122463:122432] - in_data[122495:122464];
  assign out_data[61279:61248] = in_data[122527:122496] - in_data[122559:122528];
  assign out_data[61311:61280] = in_data[122591:122560] - in_data[122623:122592];
  assign out_data[61343:61312] = in_data[122655:122624] - in_data[122687:122656];
  assign out_data[61375:61344] = in_data[122719:122688] - in_data[122751:122720];
  assign out_data[61407:61376] = in_data[122783:122752] - in_data[122815:122784];
  assign out_data[6143:6112] = in_data[12255:12224] - in_data[12287:12256];
  assign out_data[61439:61408] = in_data[122847:122816] - in_data[122879:122848];
  assign out_data[61471:61440] = in_data[122911:122880] - in_data[122943:122912];
  assign out_data[61503:61472] = in_data[122975:122944] - in_data[123007:122976];
  assign out_data[61535:61504] = in_data[123039:123008] - in_data[123071:123040];
  assign out_data[61567:61536] = in_data[123103:123072] - in_data[123135:123104];
  assign out_data[61599:61568] = in_data[123167:123136] - in_data[123199:123168];
  assign out_data[61631:61600] = in_data[123231:123200] - in_data[123263:123232];
  assign out_data[61663:61632] = in_data[123295:123264] - in_data[123327:123296];
  assign out_data[61695:61664] = in_data[123359:123328] - in_data[123391:123360];
  assign out_data[61727:61696] = in_data[123423:123392] - in_data[123455:123424];
  assign out_data[6175:6144] = in_data[12319:12288] - in_data[12351:12320];
  assign out_data[61759:61728] = in_data[123487:123456] - in_data[123519:123488];
  assign out_data[61791:61760] = in_data[123551:123520] - in_data[123583:123552];
  assign out_data[61823:61792] = in_data[123615:123584] - in_data[123647:123616];
  assign out_data[61855:61824] = in_data[123679:123648] - in_data[123711:123680];
  assign out_data[61887:61856] = in_data[123743:123712] - in_data[123775:123744];
  assign out_data[61919:61888] = in_data[123807:123776] - in_data[123839:123808];
  assign out_data[61951:61920] = in_data[123871:123840] - in_data[123903:123872];
  assign out_data[61983:61952] = in_data[123935:123904] - in_data[123967:123936];
  assign out_data[62015:61984] = in_data[123999:123968] - in_data[124031:124000];
  assign out_data[62047:62016] = in_data[124063:124032] - in_data[124095:124064];
  assign out_data[6207:6176] = in_data[12383:12352] - in_data[12415:12384];
  assign out_data[62079:62048] = in_data[124127:124096] - in_data[124159:124128];
  assign out_data[62111:62080] = in_data[124191:124160] - in_data[124223:124192];
  assign out_data[62143:62112] = in_data[124255:124224] - in_data[124287:124256];
  assign out_data[62175:62144] = in_data[124319:124288] - in_data[124351:124320];
  assign out_data[62207:62176] = in_data[124383:124352] - in_data[124415:124384];
  assign out_data[62239:62208] = in_data[124447:124416] - in_data[124479:124448];
  assign out_data[62271:62240] = in_data[124511:124480] - in_data[124543:124512];
  assign out_data[62303:62272] = in_data[124575:124544] - in_data[124607:124576];
  assign out_data[62335:62304] = in_data[124639:124608] - in_data[124671:124640];
  assign out_data[62367:62336] = in_data[124703:124672] - in_data[124735:124704];
  assign out_data[6239:6208] = in_data[12447:12416] - in_data[12479:12448];
  assign out_data[62399:62368] = in_data[124767:124736] - in_data[124799:124768];
  assign out_data[62431:62400] = in_data[124831:124800] - in_data[124863:124832];
  assign out_data[62463:62432] = in_data[124895:124864] - in_data[124927:124896];
  assign out_data[62495:62464] = in_data[124959:124928] - in_data[124991:124960];
  assign out_data[62527:62496] = in_data[125023:124992] - in_data[125055:125024];
  assign out_data[62559:62528] = in_data[125087:125056] - in_data[125119:125088];
  assign out_data[62591:62560] = in_data[125151:125120] - in_data[125183:125152];
  assign out_data[62623:62592] = in_data[125215:125184] - in_data[125247:125216];
  assign out_data[62655:62624] = in_data[125279:125248] - in_data[125311:125280];
  assign out_data[62687:62656] = in_data[125343:125312] - in_data[125375:125344];
  assign out_data[6271:6240] = in_data[12511:12480] - in_data[12543:12512];
  assign out_data[62719:62688] = in_data[125407:125376] - in_data[125439:125408];
  assign out_data[62751:62720] = in_data[125471:125440] - in_data[125503:125472];
  assign out_data[62783:62752] = in_data[125535:125504] - in_data[125567:125536];
  assign out_data[62815:62784] = in_data[125599:125568] - in_data[125631:125600];
  assign out_data[62847:62816] = in_data[125663:125632] - in_data[125695:125664];
  assign out_data[62879:62848] = in_data[125727:125696] - in_data[125759:125728];
  assign out_data[62911:62880] = in_data[125791:125760] - in_data[125823:125792];
  assign out_data[62943:62912] = in_data[125855:125824] - in_data[125887:125856];
  assign out_data[62975:62944] = in_data[125919:125888] - in_data[125951:125920];
  assign out_data[63007:62976] = in_data[125983:125952] - in_data[126015:125984];
  assign out_data[6303:6272] = in_data[12575:12544] - in_data[12607:12576];
  assign out_data[63039:63008] = in_data[126047:126016] - in_data[126079:126048];
  assign out_data[63071:63040] = in_data[126111:126080] - in_data[126143:126112];
  assign out_data[63103:63072] = in_data[126175:126144] - in_data[126207:126176];
  assign out_data[63135:63104] = in_data[126239:126208] - in_data[126271:126240];
  assign out_data[63167:63136] = in_data[126303:126272] - in_data[126335:126304];
  assign out_data[63199:63168] = in_data[126367:126336] - in_data[126399:126368];
  assign out_data[63231:63200] = in_data[126431:126400] - in_data[126463:126432];
  assign out_data[63263:63232] = in_data[126495:126464] - in_data[126527:126496];
  assign out_data[63295:63264] = in_data[126559:126528] - in_data[126591:126560];
  assign out_data[63327:63296] = in_data[126623:126592] - in_data[126655:126624];
  assign out_data[6335:6304] = in_data[12639:12608] - in_data[12671:12640];
  assign out_data[63359:63328] = in_data[126687:126656] - in_data[126719:126688];
  assign out_data[63391:63360] = in_data[126751:126720] - in_data[126783:126752];
  assign out_data[63423:63392] = in_data[126815:126784] - in_data[126847:126816];
  assign out_data[63455:63424] = in_data[126879:126848] - in_data[126911:126880];
  assign out_data[63487:63456] = in_data[126943:126912] - in_data[126975:126944];
  assign out_data[63519:63488] = in_data[127007:126976] - in_data[127039:127008];
  assign out_data[63551:63520] = in_data[127071:127040] - in_data[127103:127072];
  assign out_data[63583:63552] = in_data[127135:127104] - in_data[127167:127136];
  assign out_data[63615:63584] = in_data[127199:127168] - in_data[127231:127200];
  assign out_data[63647:63616] = in_data[127263:127232] - in_data[127295:127264];
  assign out_data[6367:6336] = in_data[12703:12672] - in_data[12735:12704];
  assign out_data[63679:63648] = in_data[127327:127296] - in_data[127359:127328];
  assign out_data[63711:63680] = in_data[127391:127360] - in_data[127423:127392];
  assign out_data[63743:63712] = in_data[127455:127424] - in_data[127487:127456];
  assign out_data[63775:63744] = in_data[127519:127488] - in_data[127551:127520];
  assign out_data[63807:63776] = in_data[127583:127552] - in_data[127615:127584];
  assign out_data[63839:63808] = in_data[127647:127616] - in_data[127679:127648];
  assign out_data[63871:63840] = in_data[127711:127680] - in_data[127743:127712];
  assign out_data[63903:63872] = in_data[127775:127744] - in_data[127807:127776];
  assign out_data[63935:63904] = in_data[127839:127808] - in_data[127871:127840];
  assign out_data[63967:63936] = in_data[127903:127872] - in_data[127935:127904];
  assign out_data[63:32] = in_data[95:64] - in_data[127:96];
  assign out_data[639:608] = in_data[1247:1216] - in_data[1279:1248];
  assign out_data[6399:6368] = in_data[12767:12736] - in_data[12799:12768];
  assign out_data[63999:63968] = in_data[127967:127936] - in_data[127999:127968];
  assign out_data[64031:64000] = in_data[128031:128000] - in_data[128063:128032];
  assign out_data[64063:64032] = in_data[128095:128064] - in_data[128127:128096];
  assign out_data[64095:64064] = in_data[128159:128128] - in_data[128191:128160];
  assign out_data[64127:64096] = in_data[128223:128192] - in_data[128255:128224];
  assign out_data[64159:64128] = in_data[128287:128256] - in_data[128319:128288];
  assign out_data[64191:64160] = in_data[128351:128320] - in_data[128383:128352];
  assign out_data[64223:64192] = in_data[128415:128384] - in_data[128447:128416];
  assign out_data[64255:64224] = in_data[128479:128448] - in_data[128511:128480];
  assign out_data[64287:64256] = in_data[128543:128512] - in_data[128575:128544];
  assign out_data[6431:6400] = in_data[12831:12800] - in_data[12863:12832];
  assign out_data[64319:64288] = in_data[128607:128576] - in_data[128639:128608];
  assign out_data[64351:64320] = in_data[128671:128640] - in_data[128703:128672];
  assign out_data[64383:64352] = in_data[128735:128704] - in_data[128767:128736];
  assign out_data[64415:64384] = in_data[128799:128768] - in_data[128831:128800];
  assign out_data[64447:64416] = in_data[128863:128832] - in_data[128895:128864];
  assign out_data[64479:64448] = in_data[128927:128896] - in_data[128959:128928];
  assign out_data[64511:64480] = in_data[128991:128960] - in_data[129023:128992];
  assign out_data[64543:64512] = in_data[129055:129024] - in_data[129087:129056];
  assign out_data[64575:64544] = in_data[129119:129088] - in_data[129151:129120];
  assign out_data[64607:64576] = in_data[129183:129152] - in_data[129215:129184];
  assign out_data[6463:6432] = in_data[12895:12864] - in_data[12927:12896];
  assign out_data[64639:64608] = in_data[129247:129216] - in_data[129279:129248];
  assign out_data[64671:64640] = in_data[129311:129280] - in_data[129343:129312];
  assign out_data[64703:64672] = in_data[129375:129344] - in_data[129407:129376];
  assign out_data[64735:64704] = in_data[129439:129408] - in_data[129471:129440];
  assign out_data[64767:64736] = in_data[129503:129472] - in_data[129535:129504];
  assign out_data[64799:64768] = in_data[129567:129536] - in_data[129599:129568];
  assign out_data[64831:64800] = in_data[129631:129600] - in_data[129663:129632];
  assign out_data[64863:64832] = in_data[129695:129664] - in_data[129727:129696];
  assign out_data[64895:64864] = in_data[129759:129728] - in_data[129791:129760];
  assign out_data[64927:64896] = in_data[129823:129792] - in_data[129855:129824];
  assign out_data[6495:6464] = in_data[12959:12928] - in_data[12991:12960];
  assign out_data[64959:64928] = in_data[129887:129856] - in_data[129919:129888];
  assign out_data[64991:64960] = in_data[129951:129920] - in_data[129983:129952];
  assign out_data[65023:64992] = in_data[130015:129984] - in_data[130047:130016];
  assign out_data[65055:65024] = in_data[130079:130048] - in_data[130111:130080];
  assign out_data[65087:65056] = in_data[130143:130112] - in_data[130175:130144];
  assign out_data[65119:65088] = in_data[130207:130176] - in_data[130239:130208];
  assign out_data[65151:65120] = in_data[130271:130240] - in_data[130303:130272];
  assign out_data[65183:65152] = in_data[130335:130304] - in_data[130367:130336];
  assign out_data[65215:65184] = in_data[130399:130368] - in_data[130431:130400];
  assign out_data[65247:65216] = in_data[130463:130432] - in_data[130495:130464];
  assign out_data[6527:6496] = in_data[13023:12992] - in_data[13055:13024];
  assign out_data[65279:65248] = in_data[130527:130496] - in_data[130559:130528];
  assign out_data[65311:65280] = in_data[130591:130560] - in_data[130623:130592];
  assign out_data[65343:65312] = in_data[130655:130624] - in_data[130687:130656];
  assign out_data[65375:65344] = in_data[130719:130688] - in_data[130751:130720];
  assign out_data[65407:65376] = in_data[130783:130752] - in_data[130815:130784];
  assign out_data[65439:65408] = in_data[130847:130816] - in_data[130879:130848];
  assign out_data[65471:65440] = in_data[130911:130880] - in_data[130943:130912];
  assign out_data[65503:65472] = in_data[130975:130944] - in_data[131007:130976];
  assign out_data[65535:65504] = in_data[131039:131008] - in_data[131071:131040];
  assign out_data[65567:65536] = in_data[131103:131072] - in_data[131135:131104];
  assign out_data[6559:6528] = in_data[13087:13056] - in_data[13119:13088];
  assign out_data[65599:65568] = in_data[131167:131136] - in_data[131199:131168];
  assign out_data[65631:65600] = in_data[131231:131200] - in_data[131263:131232];
  assign out_data[65663:65632] = in_data[131295:131264] - in_data[131327:131296];
  assign out_data[65695:65664] = in_data[131359:131328] - in_data[131391:131360];
  assign out_data[65727:65696] = in_data[131423:131392] - in_data[131455:131424];
  assign out_data[65759:65728] = in_data[131487:131456] - in_data[131519:131488];
  assign out_data[65791:65760] = in_data[131551:131520] - in_data[131583:131552];
  assign out_data[65823:65792] = in_data[131615:131584] - in_data[131647:131616];
  assign out_data[65855:65824] = in_data[131679:131648] - in_data[131711:131680];
  assign out_data[65887:65856] = in_data[131743:131712] - in_data[131775:131744];
  assign out_data[6591:6560] = in_data[13151:13120] - in_data[13183:13152];
  assign out_data[65919:65888] = in_data[131807:131776] - in_data[131839:131808];
  assign out_data[65951:65920] = in_data[131871:131840] - in_data[131903:131872];
  assign out_data[65983:65952] = in_data[131935:131904] - in_data[131967:131936];
  assign out_data[66015:65984] = in_data[131999:131968] - in_data[132031:132000];
  assign out_data[66047:66016] = in_data[132063:132032] - in_data[132095:132064];
  assign out_data[66079:66048] = in_data[132127:132096] - in_data[132159:132128];
  assign out_data[66111:66080] = in_data[132191:132160] - in_data[132223:132192];
  assign out_data[66143:66112] = in_data[132255:132224] - in_data[132287:132256];
  assign out_data[66175:66144] = in_data[132319:132288] - in_data[132351:132320];
  assign out_data[66207:66176] = in_data[132383:132352] - in_data[132415:132384];
  assign out_data[6623:6592] = in_data[13215:13184] - in_data[13247:13216];
  assign out_data[66239:66208] = in_data[132447:132416] - in_data[132479:132448];
  assign out_data[66271:66240] = in_data[132511:132480] - in_data[132543:132512];
  assign out_data[66303:66272] = in_data[132575:132544] - in_data[132607:132576];
  assign out_data[66335:66304] = in_data[132639:132608] - in_data[132671:132640];
  assign out_data[66367:66336] = in_data[132703:132672] - in_data[132735:132704];
  assign out_data[66399:66368] = in_data[132767:132736] - in_data[132799:132768];
  assign out_data[66431:66400] = in_data[132831:132800] - in_data[132863:132832];
  assign out_data[66463:66432] = in_data[132895:132864] - in_data[132927:132896];
  assign out_data[66495:66464] = in_data[132959:132928] - in_data[132991:132960];
  assign out_data[66527:66496] = in_data[133023:132992] - in_data[133055:133024];
  assign out_data[6655:6624] = in_data[13279:13248] - in_data[13311:13280];
  assign out_data[66559:66528] = in_data[133087:133056] - in_data[133119:133088];
  assign out_data[66591:66560] = in_data[133151:133120] - in_data[133183:133152];
  assign out_data[66623:66592] = in_data[133215:133184] - in_data[133247:133216];
  assign out_data[66655:66624] = in_data[133279:133248] - in_data[133311:133280];
  assign out_data[66687:66656] = in_data[133343:133312] - in_data[133375:133344];
  assign out_data[66719:66688] = in_data[133407:133376] - in_data[133439:133408];
  assign out_data[66751:66720] = in_data[133471:133440] - in_data[133503:133472];
  assign out_data[66783:66752] = in_data[133535:133504] - in_data[133567:133536];
  assign out_data[66815:66784] = in_data[133599:133568] - in_data[133631:133600];
  assign out_data[66847:66816] = in_data[133663:133632] - in_data[133695:133664];
  assign out_data[6687:6656] = in_data[13343:13312] - in_data[13375:13344];
  assign out_data[66879:66848] = in_data[133727:133696] - in_data[133759:133728];
  assign out_data[66911:66880] = in_data[133791:133760] - in_data[133823:133792];
  assign out_data[66943:66912] = in_data[133855:133824] - in_data[133887:133856];
  assign out_data[66975:66944] = in_data[133919:133888] - in_data[133951:133920];
  assign out_data[67007:66976] = in_data[133983:133952] - in_data[134015:133984];
  assign out_data[67039:67008] = in_data[134047:134016] - in_data[134079:134048];
  assign out_data[67071:67040] = in_data[134111:134080] - in_data[134143:134112];
  assign out_data[67103:67072] = in_data[134175:134144] - in_data[134207:134176];
  assign out_data[67135:67104] = in_data[134239:134208] - in_data[134271:134240];
  assign out_data[67167:67136] = in_data[134303:134272] - in_data[134335:134304];
  assign out_data[671:640] = in_data[1311:1280] - in_data[1343:1312];
  assign out_data[6719:6688] = in_data[13407:13376] - in_data[13439:13408];
  assign out_data[67199:67168] = in_data[134367:134336] - in_data[134399:134368];
  assign out_data[67231:67200] = in_data[134431:134400] - in_data[134463:134432];
  assign out_data[67263:67232] = in_data[134495:134464] - in_data[134527:134496];
  assign out_data[67295:67264] = in_data[134559:134528] - in_data[134591:134560];
  assign out_data[67327:67296] = in_data[134623:134592] - in_data[134655:134624];
  assign out_data[67359:67328] = in_data[134687:134656] - in_data[134719:134688];
  assign out_data[67391:67360] = in_data[134751:134720] - in_data[134783:134752];
  assign out_data[67423:67392] = in_data[134815:134784] - in_data[134847:134816];
  assign out_data[67455:67424] = in_data[134879:134848] - in_data[134911:134880];
  assign out_data[67487:67456] = in_data[134943:134912] - in_data[134975:134944];
  assign out_data[6751:6720] = in_data[13471:13440] - in_data[13503:13472];
  assign out_data[67519:67488] = in_data[135007:134976] - in_data[135039:135008];
  assign out_data[67551:67520] = in_data[135071:135040] - in_data[135103:135072];
  assign out_data[67583:67552] = in_data[135135:135104] - in_data[135167:135136];
  assign out_data[67615:67584] = in_data[135199:135168] - in_data[135231:135200];
  assign out_data[67647:67616] = in_data[135263:135232] - in_data[135295:135264];
  assign out_data[67679:67648] = in_data[135327:135296] - in_data[135359:135328];
  assign out_data[67711:67680] = in_data[135391:135360] - in_data[135423:135392];
  assign out_data[67743:67712] = in_data[135455:135424] - in_data[135487:135456];
  assign out_data[67775:67744] = in_data[135519:135488] - in_data[135551:135520];
  assign out_data[67807:67776] = in_data[135583:135552] - in_data[135615:135584];
  assign out_data[6783:6752] = in_data[13535:13504] - in_data[13567:13536];
  assign out_data[67839:67808] = in_data[135647:135616] - in_data[135679:135648];
  assign out_data[67871:67840] = in_data[135711:135680] - in_data[135743:135712];
  assign out_data[67903:67872] = in_data[135775:135744] - in_data[135807:135776];
  assign out_data[67935:67904] = in_data[135839:135808] - in_data[135871:135840];
  assign out_data[67967:67936] = in_data[135903:135872] - in_data[135935:135904];
  assign out_data[67999:67968] = in_data[135967:135936] - in_data[135999:135968];
  assign out_data[68031:68000] = in_data[136031:136000] - in_data[136063:136032];
  assign out_data[68063:68032] = in_data[136095:136064] - in_data[136127:136096];
  assign out_data[68095:68064] = in_data[136159:136128] - in_data[136191:136160];
  assign out_data[68127:68096] = in_data[136223:136192] - in_data[136255:136224];
  assign out_data[6815:6784] = in_data[13599:13568] - in_data[13631:13600];
  assign out_data[68159:68128] = in_data[136287:136256] - in_data[136319:136288];
  assign out_data[68191:68160] = in_data[136351:136320] - in_data[136383:136352];
  assign out_data[68223:68192] = in_data[136415:136384] - in_data[136447:136416];
  assign out_data[68255:68224] = in_data[136479:136448] - in_data[136511:136480];
  assign out_data[68287:68256] = in_data[136543:136512] - in_data[136575:136544];
  assign out_data[68319:68288] = in_data[136607:136576] - in_data[136639:136608];
  assign out_data[68351:68320] = in_data[136671:136640] - in_data[136703:136672];
  assign out_data[68383:68352] = in_data[136735:136704] - in_data[136767:136736];
  assign out_data[68415:68384] = in_data[136799:136768] - in_data[136831:136800];
  assign out_data[68447:68416] = in_data[136863:136832] - in_data[136895:136864];
  assign out_data[6847:6816] = in_data[13663:13632] - in_data[13695:13664];
  assign out_data[68479:68448] = in_data[136927:136896] - in_data[136959:136928];
  assign out_data[68511:68480] = in_data[136991:136960] - in_data[137023:136992];
  assign out_data[68543:68512] = in_data[137055:137024] - in_data[137087:137056];
  assign out_data[68575:68544] = in_data[137119:137088] - in_data[137151:137120];
  assign out_data[68607:68576] = in_data[137183:137152] - in_data[137215:137184];
  assign out_data[68639:68608] = in_data[137247:137216] - in_data[137279:137248];
  assign out_data[68671:68640] = in_data[137311:137280] - in_data[137343:137312];
  assign out_data[68703:68672] = in_data[137375:137344] - in_data[137407:137376];
  assign out_data[68735:68704] = in_data[137439:137408] - in_data[137471:137440];
  assign out_data[68767:68736] = in_data[137503:137472] - in_data[137535:137504];
  assign out_data[6879:6848] = in_data[13727:13696] - in_data[13759:13728];
  assign out_data[68799:68768] = in_data[137567:137536] - in_data[137599:137568];
  assign out_data[68831:68800] = in_data[137631:137600] - in_data[137663:137632];
  assign out_data[68863:68832] = in_data[137695:137664] - in_data[137727:137696];
  assign out_data[68895:68864] = in_data[137759:137728] - in_data[137791:137760];
  assign out_data[68927:68896] = in_data[137823:137792] - in_data[137855:137824];
  assign out_data[68959:68928] = in_data[137887:137856] - in_data[137919:137888];
  assign out_data[68991:68960] = in_data[137951:137920] - in_data[137983:137952];
  assign out_data[69023:68992] = in_data[138015:137984] - in_data[138047:138016];
  assign out_data[69055:69024] = in_data[138079:138048] - in_data[138111:138080];
  assign out_data[69087:69056] = in_data[138143:138112] - in_data[138175:138144];
  assign out_data[6911:6880] = in_data[13791:13760] - in_data[13823:13792];
  assign out_data[69119:69088] = in_data[138207:138176] - in_data[138239:138208];
  assign out_data[69151:69120] = in_data[138271:138240] - in_data[138303:138272];
  assign out_data[69183:69152] = in_data[138335:138304] - in_data[138367:138336];
  assign out_data[69215:69184] = in_data[138399:138368] - in_data[138431:138400];
  assign out_data[69247:69216] = in_data[138463:138432] - in_data[138495:138464];
  assign out_data[69279:69248] = in_data[138527:138496] - in_data[138559:138528];
  assign out_data[69311:69280] = in_data[138591:138560] - in_data[138623:138592];
  assign out_data[69343:69312] = in_data[138655:138624] - in_data[138687:138656];
  assign out_data[69375:69344] = in_data[138719:138688] - in_data[138751:138720];
  assign out_data[69407:69376] = in_data[138783:138752] - in_data[138815:138784];
  assign out_data[6943:6912] = in_data[13855:13824] - in_data[13887:13856];
  assign out_data[69439:69408] = in_data[138847:138816] - in_data[138879:138848];
  assign out_data[69471:69440] = in_data[138911:138880] - in_data[138943:138912];
  assign out_data[69503:69472] = in_data[138975:138944] - in_data[139007:138976];
  assign out_data[69535:69504] = in_data[139039:139008] - in_data[139071:139040];
  assign out_data[69567:69536] = in_data[139103:139072] - in_data[139135:139104];
  assign out_data[69599:69568] = in_data[139167:139136] - in_data[139199:139168];
  assign out_data[69631:69600] = in_data[139231:139200] - in_data[139263:139232];
  assign out_data[69663:69632] = in_data[139295:139264] - in_data[139327:139296];
  assign out_data[69695:69664] = in_data[139359:139328] - in_data[139391:139360];
  assign out_data[69727:69696] = in_data[139423:139392] - in_data[139455:139424];
  assign out_data[6975:6944] = in_data[13919:13888] - in_data[13951:13920];
  assign out_data[69759:69728] = in_data[139487:139456] - in_data[139519:139488];
  assign out_data[69791:69760] = in_data[139551:139520] - in_data[139583:139552];
  assign out_data[69823:69792] = in_data[139615:139584] - in_data[139647:139616];
  assign out_data[69855:69824] = in_data[139679:139648] - in_data[139711:139680];
  assign out_data[69887:69856] = in_data[139743:139712] - in_data[139775:139744];
  assign out_data[69919:69888] = in_data[139807:139776] - in_data[139839:139808];
  assign out_data[69951:69920] = in_data[139871:139840] - in_data[139903:139872];
  assign out_data[69983:69952] = in_data[139935:139904] - in_data[139967:139936];
  assign out_data[70015:69984] = in_data[139999:139968] - in_data[140031:140000];
  assign out_data[70047:70016] = in_data[140063:140032] - in_data[140095:140064];
  assign out_data[7007:6976] = in_data[13983:13952] - in_data[14015:13984];
  assign out_data[70079:70048] = in_data[140127:140096] - in_data[140159:140128];
  assign out_data[70111:70080] = in_data[140191:140160] - in_data[140223:140192];
  assign out_data[70143:70112] = in_data[140255:140224] - in_data[140287:140256];
  assign out_data[70175:70144] = in_data[140319:140288] - in_data[140351:140320];
  assign out_data[70207:70176] = in_data[140383:140352] - in_data[140415:140384];
  assign out_data[70239:70208] = in_data[140447:140416] - in_data[140479:140448];
  assign out_data[70271:70240] = in_data[140511:140480] - in_data[140543:140512];
  assign out_data[70303:70272] = in_data[140575:140544] - in_data[140607:140576];
  assign out_data[70335:70304] = in_data[140639:140608] - in_data[140671:140640];
  assign out_data[70367:70336] = in_data[140703:140672] - in_data[140735:140704];
  assign out_data[703:672] = in_data[1375:1344] - in_data[1407:1376];
  assign out_data[7039:7008] = in_data[14047:14016] - in_data[14079:14048];
  assign out_data[70399:70368] = in_data[140767:140736] - in_data[140799:140768];
  assign out_data[70431:70400] = in_data[140831:140800] - in_data[140863:140832];
  assign out_data[70463:70432] = in_data[140895:140864] - in_data[140927:140896];
  assign out_data[70495:70464] = in_data[140959:140928] - in_data[140991:140960];
  assign out_data[70527:70496] = in_data[141023:140992] - in_data[141055:141024];
  assign out_data[70559:70528] = in_data[141087:141056] - in_data[141119:141088];
  assign out_data[70591:70560] = in_data[141151:141120] - in_data[141183:141152];
  assign out_data[70623:70592] = in_data[141215:141184] - in_data[141247:141216];
  assign out_data[70655:70624] = in_data[141279:141248] - in_data[141311:141280];
  assign out_data[70687:70656] = in_data[141343:141312] - in_data[141375:141344];
  assign out_data[7071:7040] = in_data[14111:14080] - in_data[14143:14112];
  assign out_data[70719:70688] = in_data[141407:141376] - in_data[141439:141408];
  assign out_data[70751:70720] = in_data[141471:141440] - in_data[141503:141472];
  assign out_data[70783:70752] = in_data[141535:141504] - in_data[141567:141536];
  assign out_data[70815:70784] = in_data[141599:141568] - in_data[141631:141600];
  assign out_data[70847:70816] = in_data[141663:141632] - in_data[141695:141664];
  assign out_data[70879:70848] = in_data[141727:141696] - in_data[141759:141728];
  assign out_data[70911:70880] = in_data[141791:141760] - in_data[141823:141792];
  assign out_data[70943:70912] = in_data[141855:141824] - in_data[141887:141856];
  assign out_data[70975:70944] = in_data[141919:141888] - in_data[141951:141920];
  assign out_data[71007:70976] = in_data[141983:141952] - in_data[142015:141984];
  assign out_data[7103:7072] = in_data[14175:14144] - in_data[14207:14176];
  assign out_data[71039:71008] = in_data[142047:142016] - in_data[142079:142048];
  assign out_data[71071:71040] = in_data[142111:142080] - in_data[142143:142112];
  assign out_data[71103:71072] = in_data[142175:142144] - in_data[142207:142176];
  assign out_data[71135:71104] = in_data[142239:142208] - in_data[142271:142240];
  assign out_data[71167:71136] = in_data[142303:142272] - in_data[142335:142304];
  assign out_data[71199:71168] = in_data[142367:142336] - in_data[142399:142368];
  assign out_data[71231:71200] = in_data[142431:142400] - in_data[142463:142432];
  assign out_data[71263:71232] = in_data[142495:142464] - in_data[142527:142496];
  assign out_data[71295:71264] = in_data[142559:142528] - in_data[142591:142560];
  assign out_data[71327:71296] = in_data[142623:142592] - in_data[142655:142624];
  assign out_data[7135:7104] = in_data[14239:14208] - in_data[14271:14240];
  assign out_data[71359:71328] = in_data[142687:142656] - in_data[142719:142688];
  assign out_data[71391:71360] = in_data[142751:142720] - in_data[142783:142752];
  assign out_data[71423:71392] = in_data[142815:142784] - in_data[142847:142816];
  assign out_data[71455:71424] = in_data[142879:142848] - in_data[142911:142880];
  assign out_data[71487:71456] = in_data[142943:142912] - in_data[142975:142944];
  assign out_data[71519:71488] = in_data[143007:142976] - in_data[143039:143008];
  assign out_data[71551:71520] = in_data[143071:143040] - in_data[143103:143072];
  assign out_data[71583:71552] = in_data[143135:143104] - in_data[143167:143136];
  assign out_data[71615:71584] = in_data[143199:143168] - in_data[143231:143200];
  assign out_data[71647:71616] = in_data[143263:143232] - in_data[143295:143264];
  assign out_data[7167:7136] = in_data[14303:14272] - in_data[14335:14304];
  assign out_data[71679:71648] = in_data[143327:143296] - in_data[143359:143328];
  assign out_data[71711:71680] = in_data[143391:143360] - in_data[143423:143392];
  assign out_data[71743:71712] = in_data[143455:143424] - in_data[143487:143456];
  assign out_data[71775:71744] = in_data[143519:143488] - in_data[143551:143520];
  assign out_data[71807:71776] = in_data[143583:143552] - in_data[143615:143584];
  assign out_data[71839:71808] = in_data[143647:143616] - in_data[143679:143648];
  assign out_data[71871:71840] = in_data[143711:143680] - in_data[143743:143712];
  assign out_data[71903:71872] = in_data[143775:143744] - in_data[143807:143776];
  assign out_data[71935:71904] = in_data[143839:143808] - in_data[143871:143840];
  assign out_data[71967:71936] = in_data[143903:143872] - in_data[143935:143904];
  assign out_data[7199:7168] = in_data[14367:14336] - in_data[14399:14368];
  assign out_data[71999:71968] = in_data[143967:143936] - in_data[143999:143968];
  assign out_data[72031:72000] = in_data[144031:144000] - in_data[144063:144032];
  assign out_data[72063:72032] = in_data[144095:144064] - in_data[144127:144096];
  assign out_data[72095:72064] = in_data[144159:144128] - in_data[144191:144160];
  assign out_data[72127:72096] = in_data[144223:144192] - in_data[144255:144224];
  assign out_data[72159:72128] = in_data[144287:144256] - in_data[144319:144288];
  assign out_data[72191:72160] = in_data[144351:144320] - in_data[144383:144352];
  assign out_data[72223:72192] = in_data[144415:144384] - in_data[144447:144416];
  assign out_data[72255:72224] = in_data[144479:144448] - in_data[144511:144480];
  assign out_data[72287:72256] = in_data[144543:144512] - in_data[144575:144544];
  assign out_data[7231:7200] = in_data[14431:14400] - in_data[14463:14432];
  assign out_data[72319:72288] = in_data[144607:144576] - in_data[144639:144608];
  assign out_data[72351:72320] = in_data[144671:144640] - in_data[144703:144672];
  assign out_data[72383:72352] = in_data[144735:144704] - in_data[144767:144736];
  assign out_data[72415:72384] = in_data[144799:144768] - in_data[144831:144800];
  assign out_data[72447:72416] = in_data[144863:144832] - in_data[144895:144864];
  assign out_data[72479:72448] = in_data[144927:144896] - in_data[144959:144928];
  assign out_data[72511:72480] = in_data[144991:144960] - in_data[145023:144992];
  assign out_data[72543:72512] = in_data[145055:145024] - in_data[145087:145056];
  assign out_data[72575:72544] = in_data[145119:145088] - in_data[145151:145120];
  assign out_data[72607:72576] = in_data[145183:145152] - in_data[145215:145184];
  assign out_data[7263:7232] = in_data[14495:14464] - in_data[14527:14496];
  assign out_data[72639:72608] = in_data[145247:145216] - in_data[145279:145248];
  assign out_data[72671:72640] = in_data[145311:145280] - in_data[145343:145312];
  assign out_data[72703:72672] = in_data[145375:145344] - in_data[145407:145376];
  assign out_data[72735:72704] = in_data[145439:145408] - in_data[145471:145440];
  assign out_data[72767:72736] = in_data[145503:145472] - in_data[145535:145504];
  assign out_data[72799:72768] = in_data[145567:145536] - in_data[145599:145568];
  assign out_data[72831:72800] = in_data[145631:145600] - in_data[145663:145632];
  assign out_data[72863:72832] = in_data[145695:145664] - in_data[145727:145696];
  assign out_data[72895:72864] = in_data[145759:145728] - in_data[145791:145760];
  assign out_data[72927:72896] = in_data[145823:145792] - in_data[145855:145824];
  assign out_data[7295:7264] = in_data[14559:14528] - in_data[14591:14560];
  assign out_data[72959:72928] = in_data[145887:145856] - in_data[145919:145888];
  assign out_data[72991:72960] = in_data[145951:145920] - in_data[145983:145952];
  assign out_data[73023:72992] = in_data[146015:145984] - in_data[146047:146016];
  assign out_data[73055:73024] = in_data[146079:146048] - in_data[146111:146080];
  assign out_data[73087:73056] = in_data[146143:146112] - in_data[146175:146144];
  assign out_data[73119:73088] = in_data[146207:146176] - in_data[146239:146208];
  assign out_data[73151:73120] = in_data[146271:146240] - in_data[146303:146272];
  assign out_data[73183:73152] = in_data[146335:146304] - in_data[146367:146336];
endmodule
